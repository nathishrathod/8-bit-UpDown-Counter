���� JFIF      ��(ICC_PROFILE         mntrRGB XYZ             acsp                             ��     �-                                                   	desc   �   trXYZ  d   gXYZ  x   bXYZ  �   rTRC  �   (gTRC  �   (bTRC  �   (wtpt  �   cprt  �   <mluc          enUS   X    s R G B                                                                                XYZ       o�  8�  �XYZ       b�  ��  �XYZ       $�  �  ��para        ff  �  Y  �  
[        XYZ       ��     �-mluc          enUS        G o o g l e   I n c .   2 0 1 6�� C 


�� C		��  =" ��             	�� f 
  !1"3AQaq�246Rrt���#5STUs������B���$%EVc��b��	&CFdu'7D��´Xe��������           �� @     !1AQR�Saq��"2B�����#C�3b�$DTr���   ? �� ���JuO��%u���ߙWd�<p�βY�5�����ٝ\s�����4�e����|�:��|�~�t� ��M}�����^k�{q�S����e`y��	w���}�	�'5�b�N#`���>y6_-v��\ќ��Ij�ܢ+�2�7����T� ���ˏ�Z�����$������4�w�� �����׭�7�_C��7�v���b^��gMrmܦba����}�����t���k=AK���y+���l8��ܮ����]�co߱���)nd�{\� ܖ�wp�%̓v�[�.S>��{n��ޢ��?�}S��������;�+��G�^���6�Z���u�W!�ox�G��><;��Aj.�
za+Y�Tqm�q��fq4m�����W%.��f���&c�㣦��M8�9��Q��Ǫ�w�S��w̾���#�t����rgW�_�jW��������r���,t�wX3LŦd9WVm��9���Ā�;}���tNĮ#3v���(��[���gT� �:��|�}s�>��4�Z�2zs���m�a=k�qkGo��Ecj��{�����iy��q҃���l�isZݏ>M;�6U��T�i���;^��n���T��1^uO����ۤ�_�Ό4����S�u��#d���=����� �fwNa���KP�e�@\��ho=��+S�+�3M�~U��E3��W���� �1N�� �1_Zc~�n�2�̲���Ę����lsK�&�< o���yyV��zG�Y�')��e�ӌt���N��n[�<���#b�3�i����Dg�W��n��� �T� ��~�t-�ɋӺ��J�m�u<p��|7\ևH^V�3�_�(�w��x�t��TN�9�sZ�׵����S1��&���JuO����o��2u�f�˿��t|��E���'���JuO����o��2u�f���_�>Oi}%����}�S���]c��7�N��ߙ<1��G��-/��?U'�w�S��w�+�u�f������'�5~��<E���'�������:�3~d�|�����t|�"��K��O��%:��|�u���ߙ:�3~d�Ư�'������S���N�� �D������'[�o̞�������\���w�S��w�+�u�f������'�5~��<E���'���JuO����o��2u�f���_�>Oi}%����}�S���]c��7�N��ߙ<1��G��-/��?T� �T� ��WX�|�����7�Oj���x�K�.O�I�����J�o��2u�f���_�>Oi}%����}�T��1]c��7�N��ߙ<1��G��-/��?T� ��S��w�+�u�f������'�5~��<E���'������J�o��2u�f���_�>Oi}%����|�:��|�u���ߙ:�3~d�Ư�'������S���N�� �1]c��7�N��ߙ<1��G��-/��?T� ��S��w�+�u�f������'�5~��<E���'����uO��%u���ߙ:�3~d�Ư�'������S���N�O������'[�o̞�������\���w�)�?�;�+�u�f������'�5~��<E���'���JuO��%u���ߙ:�3~d�Ư�'������S��b�S���]c��7�N��ߙ<1��G��-/��?T� ��S��w�WX�|�����7�Oj���x�K�.O�?�;����J�o��2u�f���_�>Oi}%����|�:��}��[�o̝o��2xcW�Z_Ir~�� �1N�� �1]c��7�N��ߙ<1��G��-/��?T� ��S���;�+�u�f������'�5~��<E���'���JuO��%u���ߙ:�3~d�Ư�'������S��b�S���]c��7�N��ߙ<1��G��-/��?T� �T� ��WX�|�����7�Oj���x�K�.O�?�;�����:�3~d�|�����t|�"��K��O��%:��}��[�o̝o��2xcW�Z_Ir~�� �1N�� �D������'[�o̞�������\���w�)�?�;�+�u�f������'�5~��<E���'���JuO����o��2u�f���_�>Oi}%����|�:��}��[�o̝o��2xcW�Z_Ir~�O�T� ��WX�|�����7�Oj���x�K�.O�?�;����J�o��2��;xF�eٝU1����gL�GT� ��S��w�WU���������~�{��i�zǶ\���w�S��w�+��S<�2wS<���Ú�}?(��b?�\���w�S��w�+���f��޷�ߙi�_����-����2�5k�~�À&�x��ý�!�}~�to�-tGЕj=�Kk3l�#�s)x��8��?"�k� e}zsk�i<���T!l$�����o�.��Hͧ��$�O�6ƥŜ-��֬l8��l���ݱ��W:Zj��#<��8�^�՝4jj�&��s�}?ST�\�9����E;]���;A{KT��ruu2����"��?�+�(�����HS�]sK]�`>Ŭ{�q��wz	��Y]���U��mπ�[+g��V&9�)`=`x;�5�b�4��3��h�r���#�]g�Έ�}7hz_+3�֝앶# �74��͸�����G}�v�&����-��N@�Y=��w��_S��m���&�z���ũ��K�84�0���!=����|�{�N��h�c���v�wM�1�d�N%q`��7��o���^·S���V�_���#������"cLu��~}�r��>�b�p�d���_�ڻ]�^��g�z�Pt�j�ʮҒM�G n�=�;���+���?a�/���$t_$�<���Sk������žŽ�v/�5���t����s�_��X��lH .� ;<�}۷��E�*�1�\�/+��(�5Ӛ�s�� ��D�~Ǯ��?%I�ij�2q���]r��1��k�~e�0�&�yG�즴wLul��c� �Km�
���~����+�s��/:���aګ8�c9�󜰣kܧ�1��?L����"z)��uM;T��_9&F�]�-��"g�l����o���(q}$����;#c.1��d�0�Y�ȋ��6o=��巐yW����^��=~���,Uӏk�j� �\��7�m�$��j�C^��L�t�Z�"���j�Z\�!�li��5O� �z}�j����e�W�q�t��6\���SQ���{�`����s �{˞���V��� e֚���<�GTY��$��F9v����|A��Q�}#���;w2�w�řK���v�k~e��b�M?��3��gj�T��b9~��N�:Z�����#�skc��q(��#`<#����5I����s���6:A��g�Ut�H�^���� �����/8գb[��\矧���\�:#�I��3Ӟ���/�L^��K!xˋu{mM�n�lw=�rWk���7	��)��5r��C$97�a,�^��d��>G)_�bu�eoؖg�S���Z�t���_�X�z=�qt�#�\���RԖ�Zvm��TuOhc�nK���峏��}�ۅ��y���.����4՝�~�-f��f�M8�'�yƱ��2u�e��<��Oq�n�̝g�7��G��cu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xӍcu�d�<ɼn�xלk��'Y�M�u�Ɯk��'Y�M�u�ƽ�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��4�X�g�:�2o��5���<��y�x�d�8�?Y�N�̛��'�8�7Y�N�̛��'�8�7Y�N�̛��'�8�7Y�N�̛��'�8�7Y�N�̛�� �P]���U��S�ߏB��]?�S��1�s�� �s3u���+��@.!���������I���� �l��`�96%��c��w�-^�K���f��4�F�}� �h�	� ����c���juuگv�����wX��r����� � ��GH�*�fƆ�C^$��� k@ܒv�D.�l���Z��{�� �>Bn��$����I�m�g���x� �k��Uz����1�Խb�US� |� e��&z��bG'���
��̻���a�U?�.��5t�o���j(�6h<w=���d��{y�h�/������I�S�����jhib�=׻�H�!�nĂ�O\O�,�9�x��5;2Ք��yi��k44j����c�}�W^���i�_�3��n��ڣ����d�W��D��3��A�a��Z����߈���k�t�:t�Df�L��7��F ���_��t���y|��&����o'֩� H:���_����*6=Qތu�� /Nv�39ݟ�����oh/q�2zN֞ո��9��n�v���1*[Y��8�=�4������fq9��k��58ec��s���!jA�� �~�� �"jQ�����lv��c�O�W��/��~ҵ������!t�G}gt���j<�WT��o{�{ǈlOo�~Du�~Յ5�l�d�W�!�s�I*���W����l�sE3��r�5ڊ��"��	��S��^|�����z�:�Q�y�t*�)���=�:�:��ϕ:�p��\|��y�wt*u�8�	#�*u�ʣ���|��8I�Νq���S�)�8I��S����S�>T�$�\|��y�wt��N)�H��ʝq���S�>T�$�]�N��Tw^|��ʜS��돕:�:��ϕ:��N)�H��ʝw�GwA�^|��8I��S�>Uן*u�ʜS�����*��ϕ:��N)�H��ʝw�GwAN��S�p�=q�\|�;�>T��qNG��\|�;�>T��N)�H��t돕Gu�:��N)�H��ʝw�GwA�^|��8I��S�>U�ʝy��$z�:u�ʣ���|��8I��S��^|��8I��S����S�>T�$�\|��*��ϕ:�S�����*��ϕ:��N)�H��ʝw�Gu�ʝy��$z��N�Σ���N��S�p�=q�\|�;�)ן*qNG��\|�;�)ן*qNG�>T��;�>T�ϕ8�	#�*u�ʣ��y��$z�:u�ʣ���N�>T�$�]�N��Twt�ϕ8�	#�*u�u�:��N)�H��ʝq�t�$�\|��*��ϕ;��S�p�=w�:��Q�y�^|��8I��S����S�>T�$�\|��*���N��S�p�=w�:��Q�yN��S�p�=q�]�Q�yN��S�p�=q�\|�;�>T�ϕ8�	#�*u�ʣ���N�)�8I�Νq���S�;���$z��T����,��S�+:�L�%跉���=�n�3rd���3/|���4�j�x�]���m���WD����A�?���'^|�rܦ��oWO?Ž��v��;�O��d��j;C�x<n��&����i��+�u�?���ϕZ���3��QTMs]Y�=���7�*���Q�:u�u�w�<�̿EG�ͮ��gu.�Qr�յѯ��K�d?�/���L�_�Ɵ�X��� �)� ���]�Q���ǲ��յѯ��K�d?�'�mtk�wR���K�/�?�ߙ8�̝�QX�C�����5���k�������.j_��� )~��G��'�2w�G�N�c��O������������5���k������o̼���7�N�����l{!��?�mtk�wR���I�[=~\Կ���R���7�N�߀|��5�;��d?=?�g�S��Կ���R��=�]Կ���R�����Fe�����-�蛪/���!�<o'm� <��%1���(�Q:m<s�!�?�l�k�sR���I�[]�������Pla��ߙR�B�xx��|����C����z5��K�\?�'�mtk�sR���K�#� �����{�[i˷��w�G�N�c��o������������5��K�\?�/Ц�N�;y<p�[�p��Q��C�����5?��K�\?�'�mtk�wR���K����/�<�WL���w�G�N�c��?���������_կѱ �7�v����R�0�ohߙq���f�ƳQ?�'t��ʃ� f�F� ��7�P� ����n�� -�ڢ� )Ht��K�M9����4��|1Ճ���'�v�j��ä������v�nҹDW9O����Gg[�h�9�ܚ��n����S���I�Z��[�� �E�R��� �7G�6�O�a��tcj��V��O՟�M���!3�Z��Z�� �E�RV�F� ��?�Q����a��tcj��Xt����ڟ����~��M���!5�Z��[�� �E�RV�F� ��?�Q����c��tcj�ä�����������?jl�g�	������֦��/����7����j���S�בہ�MFxC�_�������f���H:_N]�L�j�;a�ΆYGA��x��y��:��+�}%��ohuq3E8ǫ������֧��/�� �����֧����x~���~�)c�-ۓ~c�q;o 񭗫o�2��U���r�i������������֦������7����k�����V߂�o�
��Q��d>-��n�� -jo��� ){�Z��[�ߵ��R�G�o�	շ��|��ǲV�F�����k�����~�� -�o��� )}�շ�����Bw�G�N�c���[��Z����O�����֦����][~N��'|�{��=������7����j�����kto�kS~��K�.��'V߂�j=�w[�|]�Z��Z�� ���RV�F�����k�����V߂�o�	�5�;��d>-��n�� -jo��� )?�[��Z����_ium�!:����Q��C��������7�p� ����n�� -j��� )}�շ�����Bw�G�N�c�����n�� -�o��� )y�Z��[�ߵ��R�K�o�	շ��|��ǲ� V�F� ��?�p� ����n�� -�o��� )}�շ�����Bw�G�N�c�����n�� -jo��� )?�[��Z����_h�m�!:����QX�C�������ަ���� f�F� ��?�p� ������Bum�!;��'t��ſխѹ� }�o��� ){�Z���ަ����=[~N��'|�{��=�����z7����k�����n�� -j��� )}�շ�����Bw�G�N�c��O�͎��9��0� ��F� ���؎Y�LG��?�/��Q���#n�N[yڹG�S�&S�>܎@ۖ.AW�h��c���� ���b��Qr-Q\�X޳��nnWDb<� V�F�����j�����n�� -�ڢ� )C�Ǥ������� �7G�6��������x?�6o��L� V�F� ��?�Q��իѿ�O�T_�(o�a���n��^K���S�V��O����}��&��[��z�����O�����ާ��/�7����?�5�a��tcj~��i���6o����kto�oS~��I�Z��Z�ߵE�Rh���\eu��ɩKR��k��U�%�xi�=;����$i<�i_�P�j/o�L>C�+����h�k�9��������5QLDG��_�����֦��/�� �����ަ����{�u=�S��z�iS���v�<al[~���:�M=k��N�OTf)��� խѸ� }jo��� )y�Z��[�ߵ��R�K�o�	շ��^������ǲV�F�����j�����kto�kS~��K�.��'V߂�j=�wK�|[�Z��[�ߵ��R����7����k�����V߂�o�	�5�;��d>-��n����S~��K������ަ����=[~N��'|�{��=������7����k�����n�� -jo��� )}�շ�����Bw�G�N�c����[�s���ߵ��RV�F� ��7�P� ������Bum�!;��'u��ſխѿ�M�\?�'�kto�kS~��K�.��'V߂�j=�wK�|]�Z���ަ������7����k�����V߂�o�	�5�;��d>.��n�� -jo��� )?�_��z����_h�m�!:����QX�C�������֦������7����k�����V߂�o�	�5�;��d>.��n����S~��I�Z��Z�ߵ��R�G�o�	շ��|��ǲV�F� ��7�P� ��կѿ�M�T?�/�z������G̝�Q��C�� �����֦���խѿ�M�T?�/�����[~N�����l{!�o�kto�kS~��K�������7�P� ������B�o�	�5�;��d>/��~�� -�oڡ� )x�l�l;sz���?�/�z���`�;�j=�wK�n�{��0��}@�z�k���mA,YZ�rj����F[�l͏�v�[֐�( ��7_CiѾ��|�/�ч��RY�*�̃g��7��m���<��3��[�LՌK���WP6�6�ęeu��QH٧v&H�����s�;~�^K�:^�sN�����j�Z�c��ԕ����<l���	��h8��h�5�2�8c �`��
P�9�{�0�� ���c�v#���l{A��+H���:T�+�W�� ��O��bl{���@�d��Mb�d��f�jw$hjN��ԍ��\˲u���t>ʼ�;X�<�X����k~9o/잹�Ә�&�6�X�J�����dm`����8�K!5��X��GՎ�w�&�3<�"�Q\�Gk�����vr㢹RH��9el�A(�$��7ry;�-^.�2�L|�J�1��V�v�cÞ+�k�x�WH�F���i;���d�f*�m#0v�WcZ��=�f�������[�����f��|�X�/$��O���$�IQ�o��M]2�4J�5~v�6�u`����X����;�� �8v��Gq��FÒ�t�L�M-��.�G%��,۽m��Z6���ǈ�����͆NG`WБc*�e�#�,<l�Z�����{̢s�3�1v1���jZs{��5���������0O�Z.[�&�D�W��zytu,�i�c撣mYg6� [�Aܝ�G#ϴ�J]'c�d������B�c,��ws�����d7����'�;�u�gL�\�W���Z�v]=���j�A�w�э�ۋ��&�ƸF��1��k�ն�I����nʬ-��7���~D���^���5���ՉϦq� ˏ[n��{�F]#�N��j~�s<��z�ND�9q�6���i��؃�|�юNG����zA�j9*]�2���ʆ��y�H���;a� U�6��F��@�z�Ĕ��Ê�,!̚�lL�~��w���ۿ�ozS���>�K�q���S����էSb�չ�*�����3,i�޹M1\�c1���/��]���Xk��v�?�
�y�|7��gm���-�8N�;su�c��v��$#�oc�rW�X+O?W#_%0GV�w��n�}��ک��ƙ�M�adQ�m��-��μ�=h�W����i�^K+_���f�#v;����x�u֪�M3��˧(��/K���W�=��;��F�vr=�8�7&老(JC�d��;I���'��G��O�;vzT�e�6Å��b�J[<�N�\�v#ʾ���7�s�����Z�2H�nBZ�t��ہ�Do�vy6
���n'Sɨ��Ul䄹����I�<[o��G}�MQL�������sNܾg�:Ft��F�5&�ξ����M��;���8[�r����`9-OMtO��vb�[	��������uj��?s���o̭�`B��^��q\G��ź�S4̽\o/�I�#���{�oH��r�)t>�� �ޭ� �3}e-�k霞��Ô�K����J�Y1K)�c01۽�1�<qr �&��zT�g[�G�y~��ڥf���<p�װ��e�� �>�� �,��
�R��.i裋�1������k�-��&�G���q��S�����:Aՙ����z��r;^w-Y�\N�ɿ-��k��)�N��)���?f+bo�'���̍ t��%��A^���B����AY�6fs�?T�^���N�p� �([4��d�x�:W�;�&9�Ť�#�	�A��b�������qp�Ň�����/��$G�Is{��N�]� @]!�9?���������� �����{�D���i
�q�g�%��ؖ+俫/kvcX�{5�v�$���Z>��������H��V-��������	�9�Dy��� �H_�O�{���B#�������ޱE{�{?Սvo�LS�?�Bg�o�/�����R֖)��y{e�Y���Q�����m�
�Y�t��t�O`G�  ���ѹ�6���~Rgؚ��d����~�k����G%��E���D� W��������1�>��AoQ�m?=��u���R2�����t���ak��{@��ڗ<�D�qb���u������qr��uD���`[�ߗj�����S��� �|v��j�����-S��=Q[��O��� ��O��� ��\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�\Eo�� �?�_��� �?�_�H�~����=m_?}���)�j� ���柘;PD͞�u���|��}��S1�t�l~c'r<�{���c�go�n@����ڢ�]��qy�B��Kr�z��F�������f%�q�L������x�;|@��Χ��{Xx�0cّeb�:w�eG�݇����pyHyx��i���/�K)�����/�K'���F�r�ڢ���}�έ[�n������՚WD��ީM�d���F;�K#{����8����;���E�=-��req�S�O%�#�� ^y5�)W����+�n���%@�"�#d�Jec��p�BA����~�f��M)���;�:I���M��=��k4ݘ��H�摛Kcۑ��|��;�[]�\�:F�5�p��n=����-SEB��q�:�R��8��7�?�Aw����t�� �� PS�􅿽,��
�z�MS{?��]����?��Ӷ���ү��j��s�}R�~��+)�V1�x�f��'n��y�e�4WA������\�U��W�Yٌl�$�@}[k@碣�����v!,��\�<	�]#8���7q�o�|���Y��D�=^���ަ�Q4�O������z?�go	f<�"Z���c��.رǑ o��v5�C�3���w'���͚���d��^�Ѵ��s��܆���֝�� ��_!����"Y���w�au���T� ��N��T� ��\���V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� ��V���S��� �:��S��� �Ńs�B���O��� �fa,�7p��s\�=��A�i�� ��ϒ�����F�l�JpձY���$��b[ֹ�#�3o���0���O{��|�/�gC�û��6<1��O�˟��S1aI���m{��|1b䊤�6#���p���ov���Z�;A����+�
y,�<k�I�)�k�~�i�Ʉ�� ���&9�	�
�f��H"on�m�ݛ�*��Ѯ��8#t@�720�� U���Wz��;��l�Xǹ��վ#�{���	 ��♽�{ ;��Lu]�<1c�U�O��a��ќ}�w �Ƿb�(���\�GB�nc��[G�i�UP�(W|O��x��[�Af��r忍Zj�1�$Eq��GL�;��wc,2Y���T^����#{�ݷ>%��0�K����Z3��z���wѵ�NnFF�܃��e�M'�7:�t{�w�v�Gb�=�1�!sbqtm1��|��%U�*�s��M�ש�cǉ�m�呻��#n�|Hp;�����3֠ۏ�(��Y���X����Dv��q.�=�������/�Y�o�.���[y<�a�M�._s17���r��I�ʶ��_�b�V�ޖ��C+f�.̞�ۂ����׉'ꋃ�?��$�ϟ,8S��"�43ڦ��a!�,qa;l�^o�.��e.	�*��1�ucg�)�̪N���X�408���G`�n�2EV�&*�:ba|@b��uy'|%�݁�s���c޷�n�ڤht�F��`�#�����f�u��6���܃�-�غ{�ܐ�o��lG̣�G����V�^���ҽ�n�Iq�� �7Q5[�(1_�M9c�Cb\u���j�B^���x�ż���ͽ�=:��ZY����lO�5�E�	v͕��rC�-�Fv)���guN�x����r�F���a(���]� 48D7�v�޷�F+�h�~���gi�+�"������H���ϑ[�ՍK�	��F��0�@b��`au��O7pWq�n\ �Æ�^��*u����܆Þ�E�jS4�Jp=��C�r$��s�޷�JqW�Mӽ)G�rB�\�����6i$i܇��x{F��p���,x� ��L ��ܝ�w;�>U�в�bg�c�U.7��$ޑ��싍�=�7�}`�gY��mO̳��v���3�mO�3�5`���4�'����|6���3��^w<?�o̝����"0�����	�G���Os��&��+��L��*���~p��c�m�§�a�>e�s��6�ȅFX�~p�3��^w4?�o̝����"U�Y���:�Ƿ�T�<?�g̝���� �����N�?�ߝS����2���~d���6���G���;����N��l��W�G���]�oΨ�xϙxv�m��W�G���]�oέ�!�n��2������P+��m�Ӯ���Tw<?�g̽�hϙH�����N�?�ߝSܰ�	�2w,?�ĝ��?�ߝ:��~uOr��&|�ܰ�	�2
���~t��m��=����'r��&|�*��m�Ӯ���T�,?�g̝���� �����N�?�ߝSܰ�	�2w,?�ĝ��?�ߝ:��~uOr��&|�ܰ�	�2
���~t��m��=����'r��&|�*��m�Ӯ���T�,?�g̝���� ��g�oνk��� �2�Ջ�>eMf5��4����"-{���)~�TG���O_�"�׿J?#��WC�^[���r �.k=�*u��6����k�8|�Uw<^8�� �����N�?�ߜ*;����N��l��U�G�������{��~e�sC�&|Ȁ�φߝ:�|6��ܰ�	�2w,?�ğ�c�m�ӭg�oμ�Xϙ;��3�D���m�Ӯ���T�,?�g̝���� �����N�?�ߝSܰ�	�2w,?�ĝ��?�ߝ:��~uOr��&|�ܰ�	�2
���~t��m��=����'r��&|�*��m�Ӯ���T�,?�g̝���� �����N�?�ߝSܰ�	�2w,?�ĝ��?�ߝ:��~uOr��&|�ܰ�	�2
���~t��m��=����'r��&|�*��m�Ӯ���T�,?�g̝���� �����N�?�ߝSܰ�	�2w,?�ĝ��?�ߝ:��~uOr��&|�ܰ�	�2
���~t��m��=����'r��&|�*��m�Ӯ���T�,?�g̝���� �����N�?�ߝSܰ�	�2w,?�ĝ�pwa�s���,����-�Ca �'����g}��8��1㧽��>K���3��t�u��(�L+����xZh"����Ѵ��Ob�K�
Co2�5M3�V�w�r���*+����I��.�t�^�\���{m�{7[>���ٝ�L<Η�mk���k�=��sv�s�q�}�`�!^n��q
E��7�� �q�"񉒲,�Fw�¹��ېv����j�i>��}��A<�7X��29��R���a�}�y.ѱ�{�g%�z���8{�i�^�����}�Z�q��]+�Z-m� do�m�<~#���k�M���ǖ�#z��3�P�Ø�`�m��t�˱6Yq'�mϽ�/�O��vH�7^5쌥�K���|K]b�snܻ��z��W5b�-W�Rub�^���؞Oi�Bvm��.���?�8����rᴺ3��?FZ��5f���k?�&���1q8���|�ѐא���ܱ]�km�� �{�g&�����!��q�y¯��Ï)rJx��i����}��6��O�uf7��ĉ��G�S��� [�q��$���d�k�������i'�;<K�l��vc�ÏT~	�b)�;8%�F�{�C@�H/Qe�r�9��"DD@\o1�I�#���{�oH��[�}���z�����'}b��}���z�����'z�I�3�*��Wg����Dn����[�S��<16b�v�� y��#�L���G%j�톆m����#ű��o�n;T#N?z��mwD�����qp�'m��m�.Ŷ�#����R'+��/GX����*�ۄ�RY"d�0�=� s����m̍����`"�j(,�kE�l&��d�{L��w�������\>͹���D�}��U/6��uK8�!�.��A<�H�6 ���f��9�p|P9���u��[�@kfa�s�L�ъ��}���x�۞��Sb����(��?/Ey�k���naߓ��t��E�U�t�{�\ֲ0�睃�4�]��;eͯ4�sbbe�Y�*�%QV	ga 8��1���~�Bӭ}����ֈd��Գ��ckga�k\��[a㓁������}};^�긘�\��P�nR�����k����'��^h�r�S��3Sbf�Ӳ��a��,ת�ΜE��=�Z�K� ��qs�6[��aк�Q`!�]�X��+N����gXZ��˚Kv#v�w�櫋�<��%,v�}Ve�lp� ���㗋�8� ZH'm� z�ܧ���2�-���#�1��-�:���&���r��!�c�����SͶe����r��In0=�|�;w�-1��8���ƶ1F7 �y�����F꫸���Աv
b���U�	���X$��nK��u�#�� � X\�q�9�23����/NA��/�3�jǑ8��l%��g%� �Im�^�4T4q��Y�3$���z�M3�/ͼLa{:����4p�$*�Ð����j�����(�G�ٸ�Z�w�yrXK8�y���>G#�O{uns)�y�V��C���KS�~�tDv�FѻO!��c�c��y��K�x��pzCKI��M���QcOG��Ϯ%6lM4�lYx����9�� h$]�r8�"qy;T-[{�C��H9�{�h��v�"�)�/'��N���OK��G4u���'r�����8x�]����R��L�Va���p˵-��s��s��1��뚞�s���co!p��W3X��u�\�N�w��@��޺ ܆r�IH���}�Z�Okw��-KqԞc�A^VD\Zx$sC$��p%��B٠�����Ϸr�����KRe����7�P�X׮��\��!�ع� ���Eޢ�p����p����D@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKyp��$�K�}���n��Pb���g�Xws���׊͡�#��w7��l>e�����䢨ظ����޵����4�s������i��٪kɑ��\�[�6�����8��yx�]��O��|g�g� ���,�?����̄�J��8an�v5��.�/*ʺ��ᆔ�Ns-���eb�Z�l��+�{۾��qk���g�0VG�\^+):�����Q�W48���� O ]��U��,E<|-%�F��|n>RN�9P0�3�Y��V�k����G�YLr�Z��zC��C��̻ʲ�����ͥ�US<���ε�������XT��K�^�4�r�q;7���'����3��bi�ZN�����#��H��$�������nK�F�T����ŉrm�(V{]��q	/��߈q{C�;
�Qz1�śS���3��`��x�>͂i��v�{K�%�i�}	_,�W����=ď) �B�p�:�!����|�"�1���Ő9��l��Ewk�)�9�cE�j��Xò�:׀Z�NÅ���^���s���5�khl��9Z��U�.2x�N�¼н������.������+��栫g��+8A/keu�����G5Jo]�b7V�V�3��~����Zʬ�XZ頉�<�ކ��~]�凕�=�U����&���Gk�����W��J�k�S�EI�*�q����/�㌀�6�c����ܷ1�NQj���U�hv}�kI��ԗ�>�O�7Ma/�'~@o����\�n�3��m�sd)I3��ӶH�J[Ո�\�Cn�ݶ-��#%W[�̷�;��Mǯy�83����9�q�u�p��*���Q;�G�}�~9zU�f��9�o�;��� Aii�Ug�5
��n>I�C��)7-y�� ��]���<��k��lO�4�2=�dnv�x��)�~��ΜB/Y��(�2�����/�)C����q۾1�A������Y�<�]�ozvp����gk��2jl�b(�Ռ�[�Ϲ�vW�9�܉,.���5�_C�����б�u��qO��/��e��Z�Ț��G�s��*�{�8��_�_�jc;��������m����T�yz���7������^|xf�R�Q-F�ח����7�!�y�>к����nRI$��WdN�Wq=�4I�nN���]uW4�N"��LSS9I�"�b""" """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�V�[P�t��X�^���k��-�m'�r���VNXau+�f'-K"�2
��B�{7��Vݙ�㒛��w<�(�MQ�ݧuN�Ê�q��XL�|=We��=��įjΑ4��5�o$�N�8������47�O �r��#��r��g�eE��zh��~q��1?����#�R��dݭ#����9o��W��d��RЯ���ZS_��k&�lHq- v;o���O��YG�47TZ��'麵2֥ɱ�b��q�S�Uֱ����v�����ח:S��5$x�Ǖ{�����ڰ�n��i ��.j"���<[~�m���3�����e�B2m�ڦ���� � �.|���{,��)i���M?^2ѹ�0�n&�����K����<�xu�=�G��"�m�ū龓tޮ�Ϗ��b�r��6���h;4��<�i!j����tn��	%�~�ҹ�:�$��lz�̍�ܔ�j��݈抯ۢ���N��T�+Z����ϊ���������on�ol�j�b4Ɯ��|q-��p���Ҳ1�4���\��Gj�Q3�Zn�Ns=:._�:p�e5S��V�V,��uHǁ+X홻��>M�� ���E�Z���D訿���T���n``=���n|{lAV�U�8�R�E��1SzE�\�F����O���.J�!�E#��7s8Cx��Ǒ �|L�Oc�����)cr�Ƶ�s������x��C�;{vp��O�q���K��������7p�s�]��t���p4㗏e�b��3x���؎�;E4Gv�����4UO9��E\����{�oH��vE����>�Uh�xϽ�?4�PUS�?��YT�>����=AUO����e$���i�`N��ϒ�?��Z(4�%��S�u��i�^X�Lݛ.�l<�5��H>E�҆������x�0�l��m��!���"��8g���\&�fvK��&F��%k�vs��h�;	��Y%xK�x �<��U�f2�E3���.;�\���.U�薜� I����h��ټ��K���&ff��C��6OC0�a����c��H����wݻ�9/�R&���&�S�7��W�Kڵ�Z�we�VAF'�H�J[�����G0�i�L�i��M�s3M�GI=%�5n�גO��O��-V��	�#|�6��I��p<[m�>B��B�+�մ(�M���٣jI��s>Y�#�o�k~��ﺎ[����4��R_8�d⻡�	��7���	-�ý�9�)�5���?3���6�Bj��FKc�^��pf���<�����r`t���龍5Nc_����j�]Y��VD�0p�n�/�Y߲%�u�հڗ�
]��C%�nY]�o���F��ٽ��5�kk�.GR[�Ԭ�o-X8J�U��c��ӆö#v�qs�Z<���W��ٜ5j���g���!�H��L]�8��ם���.Wr�R[����lX�>�83+��Z<A�k^<�\s[�����H*�v��qYٙ[KF�-O(K$s��< ���=�+��1�zA��i��b	�)#�b�\�N�09���sce����N8�M&66���a��3��>o��֥�����3PԒ:��~�~T�f+�P�H�[U�'�]����:�MCC#��\�ҧONd�����=��
����E�i�۟x6#��:\�vtͼ�7^0�^�n�N��t�kb귌u��sZ|G��ڭj�tΚ��瞾JH3�V�Q�����#��q7�;� 8��$�G"��*��G���g7�YŰ�.5��w!k�܆m��0��m�tP� �`�L�ߏ�m.q�6�d�.�s@i�\�/<6Y+�/vN���n]�ri{��Ė���N0�e�Ud�����H�6�����9��G�kO�)q�>[3��3�u��l�C�|M��1xI�o�XxT.��X�ŷ9n�1V�j��E^/�,���\N�-u���v;���NZaak9���f��w\i�c�1X�N�v�>�z���ŇD����e�h�#p8��lvFޑu��t�c���3�|�lXwE]N��[9�s�̆����䫚k�]U��i����_Q��Ǘ��h�R<|�z�d|bA,nf�Dl�H��'��#�/W6�Ȳ�Q�c{�I_]�m#:Ʒ���	���Y��X�:���q3���׭$�=���F�;`7%�l2@A=Y�EZM7_+X־^�7����v_6�rM��j�k.ehֺ��w��<w4F9����bw��q��4���s�Z���8�yA��|M1��hپ�-���#�$��t��ܸ��1��kV��3�$�k�\�c�y�i�9�m�;���f񚷮Ը�t������dLmw���ӳ�	c�[���=�+����Zk5^�՚{$�#gBfu�4o�@Y#7��;��ñ�[�9����D@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o��P:���-��&��y��3��HO&��q|Jx�(G�+lU�)�&hp���;�H�$��vs<�lx�͙�r�JYǐ�:7U��rD�!��飅폱����~�ܕ9�x����ul��%q�JY#[j���<	Ga'�گL����˛�&���V1r�:��q����,-t2�Hn�n���r�7<�f��Pi�K,P�K�� �n�8��7��s�m��vr����{�H蹰0U���&�b��F`�	���D��+:JƓ��C��Ш�m��Z�ɡc�#ct`���\���e-SΪ3��c0�tgL:�V�'<:k�Hӳb���� ����;g9ۓ� 7����˃����|�1���T���e�
��M������>!�c���Y�橆=?�H*�d�^0m5����������M)�-�㊭��τq$Ԋ&:w� mڕ\����Cv���5�KY=������,�R����Ձ�8�`߈���xH�o����o�7�R�9�r��4!�2����!��laĆpMx�[��SL�pM&/,R��D�B�(c�ݍ�Ѹ�<������9���c�m�M��3�}s�'���gs����x�q�?8F%�^��j�2-�b�E���َ7G����ֹ�;��	�cȍ��dk��<V��ƥ�+y>�U���A�g�\F�c{6S��>FR������s��z��[�����a��^Y��8��K�����:���\X	��<<Gι��MU���j�f0�1&j+Z�8mRƌ]��C^8����l�d�y<;;� ������R��l��fN��eJy�F)&�W���Y�4��=�@K]��@<'�[H�����nu��7k��������:����{	Zxt�<u*�N)Y�c�����Y4X��[ˉ����o�m5�m �8��x� ��^հ����ÿ.:��n\��y�t1�;�ӳ�%��)kyy��^9
�����"�[��K�o��ݼ�9E�s��x�Dd�W!nIO��"�6�mn�͉t� o��7�l�Kz�8/GS���*e�"���+�+"l�ᇞ����pV� �4�S�]R���Y���' �i���=����|�m���c�?�WOпSڦgG��X�1�]#��[7�w�����&#����㕎k�#C���A���X��U�XO���1�[����)R��0�39���2�G� �c^�����fA|A��I$�� s$�"�i�@��" """ """ ""5|�YZw�K����W�~�����}��8��1�KE�� G�𙚭�J�8�Z{Xx�i�y�'D���n'=��ɹ�3�[� � r[V�����,_P)�\�)��&3j���1�ޮ]��'>�K��X#��jyg����. w.ҵ>��:�]�i�n�($�f���r̂X�$p=���@;�H+���kE�����X�������&���s�,��mX���еұ��dR4�}�s-���䴽kO'��Vc����6kMЯ;e��X�,pxgs'���n�����i,6_#[!wN����4-t��W�Zӫ��5�'5z
wqD�pY���������G���!�L�f�"5�0���;�?s�sۚ��'G�?��<d�h�3N�k���.k������ym�侓�x�QN��g1��(�15K�l��0�l^���c�v��W���&�=�c��9��\y �t7B��=�k׿F��rs�+�ݘ=�C��Osm�Y�l|\�5�Y�p�柗f&�2����y߶�]�`����)�th)��s�tp���N����8�b00U�3^K��}i{K{�q�{�v�9r�Et��β�t�k5��3!{�Y�|��6!�,F��<L'n�^@��E�:�����QU�g3��f��}��O��Ԧ���s�+dc����wؐw�*5z�_������p�U����[���6;Q�B8O.��}��v��泋���-*�SW����[=k�F��k��Ü�h�o!l�����w�����=j�_D�1��A�8�.[��y��̯9��<��!܈��K�"�u5r��46�<���S㲸��A}Gs%+f�,���qy;�����r��C:�����e3C��e�Z�-��W�>&J7�p-;�aߵ}0�gU\׾��kss2��^���;��KL�nA�.[x�8{�������p�� �ͷ滇Gx��/DajgMs���[h�`l|~> 0eE���\�7����[�ϖ����>�]�q�ǹ&��[�}���z�����'zʧ�����
�~���(1'����G�]��?ҭ�4� p_���Ď���X��"�d{cϴ�<�mUNա��Թƅ�߻5�o9�J��sx����7�p'`@ ����;	��}����i�tg��Fgt݉_=<��&�� ��>W��ɰ���0%��v�����3��+�D����h��ɤ�K4�kv���;v�L�L�8â�5LL���O�U��>�m4ح:L�mX���*�427��+;��x�ظy�U��w��rkҳZs� 26�� ���H�}�\�If��ލ4�j��*^vdտ<�d�8�d��6�o~۟*t��ָ-a���d��_q�o�Q%��A(�#�N&�}��w���ڭ��rf<�U\�ɘo�@[ҹLĘ�ы��b� p�Y�1Y��=�M�-�%�'˶�l�c����&t����4���>#Y��+�؞[�v=�`��7���Z1XyzY�A�Xfm�u�I�f���$�\{2v�<��qlQ`�.���c2�Z�N�nV��<����f�n���q۽k�i[qp<�Z.OA�4���5��B"�l�J��x�f�����!�#���q�JΗ�-�2r��\�s�D�ws��u�p�Ƿy��۝�j̦���][�]�S�:Z:1IZ��\�������ўG}���
2�D�P�zk[?iװ	25o�`��<N�a>���5���k��ք�
��8k1��fU�� ����o9+V�s1���=�3X�!%[f��?Q�,���w4n����ݷkw v�'1��ܥ�mrݚ��b�q��Nq헪<����#�c�o-�j��s��e�U��WOÅ���%�c�@$n]��rL�g5x��U����r<���5�2�xxD�Bv�\@jm�u3"�K킓��b`�<��!"㮆[��qk��@;��V�NA����fm�{/h�r�1�l�`����� �r�-S�.�C�o^nr�*7�Xܵ�L���g�$O��<�� �<��<z>���e�З#wQ��X��٣��%�$-c����<���!�S:�Q�+=��|�2��@�>(����p�H =��y�t/����Ah|��b�j�.��.ݖԆ�o�_e�X�'� c;y�w[Z[R�{ԲYZ�4�S��VZ7=�d�L�����}�#~�K����ln7��1a���+]��٢!�7�oc�-�$� b�J��-D�������s=�/ԲYX��>��Q�kI_�]�yL����MU�[f�B#kcv�s'�<�-����Y��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A�V����su�Y��g���iߑ ����G�ؖ���Y�ա�	��fB_a�������|[�c��2�Lۍе�����0�c�{�4�=��pq�2;�~�:;�����3]� �M�$���4�ذ�w� �y�H�\ִ]��Pڋ�[�R�tO�u�2��!�W���q󻸫�J����|��w� ���3���ZkL`t�gb�v�7n[6^�F�B�%���<A·\H�v#�;/Hڊ}5���͆��h%�Թ��f��ql\;�[����f:^���T~�G-G-�kg�-z���9��������ܹTbܻTrF]�ڳ?7H5����v&
wk]t�5̍�L14 �<�ݛ�tE�2G�nQ����Fsv4m`���&�~��$�wZ�^��DW�`�,���dw:��E4q=�<��+H�ߟf�GV����B<&>��hghb�l�,l���\F�v�i�|{v��L\���&���Ft�Ѿ����ݜ �ɍ�U�Cbk��M;R��5�?�l�\�?���~��`�Rd�q���2���eh�!�rӘ���7�48��8��5$�J�:�l�r�_^֟�o��z��5�����Wʸ����}�H���N��mW�[��\^I ��G[Ec���a�rZ������MN��e���ѻ�L�A޸o�;F���S��<a���I�5�dN�q;]�q%`c%�V��fţ�
C-�}��֕���d.���J��رf�}�͚����|���䁹]�N埖�н<Pג�M�G�v!��� �[s�A�,}�Y����Z��[�(:�L���"wq0����-��czӶ����t�z+��c�8c����u��L�臮�{��v� ����ĺ�;�PrW���-Y��8�<�Z�'�I�ԢZB'>H���D��і�[�m���x���/k9e.�e�eNm�;��d�e�Ts8v��dnǏn�8A�oD>���{��PV�CV�,&9�AnI��jId��Q46��3�Ǒ'�K��-E�,�����cu5ܭl}�LP�$�K`T�7�� ���q����ޡ��4�����K9
�&�ڎ)h����0w;���cs���۴��z�@7Bi�^�z�)-���f��l������N�{F�-����5�UBŋ8K��ge�i`o2�:9#�i�;���l�U"��NA�" """ """ ""5|�YZw�K����W�~�����}��8��1�N�{�X��Y�kN���|�/�οe�FZs?�:(�]���򚮦"䍙��u_��M���`�<~e�~3�MQ��D�i|E\=--�䳈���<qIU��7���K[�FG�rG=7#Ӿ��5�w]�`�O��T�U�6`��=���E�N�q�#����^��e�V��!u?E8��tncuEY,j�^���m�}i�#$��Ę�\F�7`9�%�Ct��'�ئ�,�+�ex��� r}	�9��9\�!�.܇s�A�'`^nW�:_�պ��͙Ӻm��շf<�nh����V{! �̈́ ��ǊV�ř�?�MQ���\-��n��C�Ԣ*��D��Z�pq���q���m����������R��}��4��E��MǶQ?�Q���0[ۃs� u{�;w\?���J�4��ˎ�X�N�X�m��u��@,� �q��ݏ.�q�xW����g_��G-����,m���coK3GK��L�c�~��e� ��£�V{X�p�Y�����Xv�:��bx�~�tr9�7v��}���>�p�_e���k�(�sZ~{w�Qd�:��b���j�D��$��hi� _Nt������:��[���q��ܩR٣꣑��s�fݾ$M�{�oH��vE����>�A��{j~i�����I޲��}���z�����'z�I�3�*��v���g�U�x�śy�lPegAdt�O�7wo�Oz9�7��[eQ�h~(�(*x�c�C�#��=��$� �  ��=W��|A�AYn���V���a87�Un��ޯ��-�v"�V&��4�c �@ �`����э̯p1ǈ�6��|��k I��� ^uaU�n�X���E�exc��wlL�yx����8S�/w�n��k��6�[:����qp���7W�t 6���#������|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*����G�Ef���lU��黣~��$4��`	ϕJ��j�����CY�1�ke��k�'b��6���A�c6g۳���)�F�l�x��0O��)#؃V���?��V�P֊�cf&C�kx�.;q8Gnݽ���ɂ�-��_<X��6g��c������;�02"<��+��cSi�h��ѵ`\�`��]X#��n�#~����;V���+�����Q��������#�����lA� �Ds��m��ьFjæ�b3V:/Bh�;���܋�[���/a/�Ğ�oނN�~՗��h!��T�3��r�2W�aō���(�'� {�辉5oE�'���b���Ē�d�Ӱ�p�\=�߬q�ض��8ԹlVz����������HX|��\W�7Hcqu.A�n!��-f#<�i1�[��U����>�cDF7q4�n[�n�F}��d�5���H-��%���!s߷�v���Vˎ�0	Ꮄ��_����v���z��z5n#�#�N��y��������a�c{���m��.7�Y��4f��J9p�0t�u��gk���f��{�ָl9��ʧ!�X�t��s��ny.Ђ��V{����8�!}� �����DZ��DڃM�}����᳋�����.lrO�1��tNe����۞���gz���DYlM23tV��nZ�g���B��:{�B��X�Y�4��Ė��ج�ʴ�Ev1��^U�T�Fgr[h"W�a��������������ryL�>i��ኛ��G~���J��#���������" """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���m�;V�X����
�sw�
�FL.U�n(->���wM�@n㓀$n9�*�*6ɉ���q�0�|�Z��������N:F&�l]k&yq&�;�� w�;�G�ݘvXѦr�gT��:������ͺǋOi1ϡ#�RJ'}f�h���yoۃ��Q��_�cͦIR���wDL������wy.��xsI p�F�b��NgX���W�_�N�+��u��9<�I�b9�=�������&���bq�-L�2I���=�s��	܂I'�R�Ib�ib��[����Y�!iixټ�ZH��V�'��VkS�j:�-^�k6Exk���9͐��	X{����1��I��J�o�-
��1�Mֵ����$������vﻀ� �nI4�-�だK�Q���"Y����O%�^���5y��R+�W��놘�!�Rӷ"�����Zf7�<Drу3(��K�Z6>1�ZI�W�9���ֵ�1���粧Qt����.���a҈��[�F�n�p�y�}��o̖��naѽ����֎-�߀�̡�a4���3sb��e� m�*8۳g���G?��,�Ij]��d�V���s�xc�]���8m����J����L�b�OC4����!W+�\��8862_����΂i�4��'.�4�P��7Ma�m��m�ef�Jc�l5qx��6qi���Z��7�@}�߷�k��S�b�mׯ��yٓ�ڤ������H�/%_�tрԗ����m[�nw��	�A#��6Bݸ^"Oh�~H5�+��Ӻ�-��=�Ak �U����DŭkcǍ�<O�wz9�]>��|t�e�5��']a�C�e~�q8��� �����a�tI,�f��,�%
��h��Z����4m��w��S������έJ����e��g�����w���h6�f�~���٪_�� �� �#a�����S>��b{5K�������R�7���,���|��3���'�T�� i�	��/����1�`|�Z�k�^͚�c�� AX���`�@������9�ث\��&���ĹcܓzG��Rw��auwIY�toۉ�~÷-����rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���h�����g�U��B�6mϐ�'|�k�1�9�;?�M�����øo-���}������Y��h���q��b�ø�qp��v���m�>ݷJ���R
���_0k��5�3Mݎ����bq�/��G26�%a�Y#��#�8�xI��y/��b�U34'�z�V����L��H��<�A��6���vK!j+��b�Ϲ�X��&u�	C^Z$.ؑ����d$��O��,l�[�K8�%��s��[d堷a���������7�2b>�Z�W�__þ����>e����5�*�f�Bၶ寊��R��6I8��s_ɻ��$s/��*,��+�2r��9�Uc�ƈ�Df}�;p�i*4����M��X�Rt��u.�n�k�u���aia�v��?nL���!ð�7t�S�3Zv�H��4Xl �Pc�۫���������T���N���.�c�}�C���p�.Xq"'Ih��#��(����Jhh�Pjl�u���b7�͎g���dOp;�ӿ�}�kZnS76��ϖvX6C�k���L�w3#�ޯs)~�n��l�mO��V�qvt��&z�qbH�ց�C��t�n��<�$�;�������G3���"��F�-���=����6�|\����Y��A~��=�UY��B�͡)���b����#��W�5nt�����m�I��v����"1����;qù���1�����пJ��g�<Nr�B͹q���ZR[n����nx�I�`ynH o�\�Y�M[Ђ��F����A�Q�x��3+M���ve�%��6�aӺ�v���<r���=��H���nV���t�gDj�I'lT���;���i������ُ���}����w�"?�n�j�ջ�����;���w��s�Ը��Ԛ���x�Pf&}��
\t�k9�E��6���ѳgi<[?p6܎�[�^p ��Ce5ޫ�O����{U�E�ٛR�%fI�l��ٶ�ۮ!�<%�;�ۨ�\S�NV'(,W�c˶f�͍�{>��7o�����^������"!MΨ���ǳ� H7�o1w�l��T�����qi�;�V�V#�DVD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�ZƬ�[�ݫp�b}�gG����O/�ʅ�sc �9rt�f8�xs�}���	�[��ð��?�R'�Gcu���,g� ��	� �:\Ԓi�3^�3Ӌ|�H�e����c\C۳���w���|�J��vs&�b�M����� y�QlVa��#���;��.��u,�*��.~L|4��Z������`��?:�����H��#��E�K l���i'���۷�mL�G8�z*�#�9q�gO9�XN�1b��LT�ʌ~���,�w����p��un��R���̶K�~#��7Qc�wi�ұ��k:N"l�<�kdЙM���p�\�2�Þ�_4e��4����� ���q�
���雘�CBL\�-���Wtn�g4� ��N�� �i5S�֓U��q�I-
�hlH��k��y۵�s����_:j���)����Q��I����\{����d�2&�q7���]�o��.��{���L~ټl-��R�����#~|� �{v*5���j�+�1y*�U���5[��kc�G#^�=�y��11��11(ގ5��U�Ԙ�Rм�[���8��A(�>3�s��x��=�aش~�zC�b��P����_Zۤ��,Z2X,-��{CKC7'go�õo��79��_g���P����\��29�]���rq���������|2��R�)�2?�oi,�s�;��;s�v}�>�P�Ө�f$�"㠓#��;�3V9$Jz͋d��5�u�;�	��"uN��:x�Ui��S��lG)gs��H$H��{��l;>�n"�t�dS�,J�	&����	�r=*f��b�Jd���{������ihr��3��9���m.$٧ӭ~,��I0n��D�H��p�v������i��cZ���[X�22�������doهn'x_�:΃�4ڑ�&N�xJ�7�#2���F�	xg}���*Uߧ9��QG�sU��D�����Y,e��`G#� �3����6�g'OU��{��cC�@��G5�h�>ٱ>�E��N��sE��K��>?��o�[�ek��*V���8V�,A7u��,NsZױ���IA�{G�)�,�K;��d/�lUz�KN�U4��C]��m��ŷ5��3,D�#sd��9�i�8���D@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ٱ|l�a&k#c�gn�07�Ej=1���K�"���h`229�	!�h����bӜ��3�}@�M����-���]|��F�2>}��o#���D���G'�r"���͈�!#^ȡE�l9���;7q������k_t-�%bYߵ�����7u��[e}K��NŸ2�f�^1,��a�dL-�s��ݝ��s^��x��,��R��� ��,1� F�c����ăP��R�{Qd�wN6�*Y%t��`��7ۑ<���f[Hi��,�K��IdE�}���6��-;w�p��<cu�c�T���F�7*�7�z�	�ܜ9{�#�К��Gv��08��ei����n����ɲbM+�vJ�衽Zj�G l�l�ǿ^ ���X�t��N�Y*]0�l��&�I<s������x��_Rb-����R���X�a������o�5& �e!��n>W@���:�#Z��k�#�����WԽ�խI,��xl���G���7sA�srVt>�K��e%�g lMa��$����ٹs����6pۚ�0e�ڿf�7+�v�i��r��E�7oAݻ�c~�}�k\�G���#�e��22c�u���wx��#x{6���H�x�	�ҘlM��23٢e�d����#Z�˘١lX��34d��k�Q�s��8O��y)I9�����w���Mbi�^�9*����)�t��1"��͍��Ee�=�L�1���C\�2��� ����ۅ��Ă7<��n��6D�FV |� �w�^�/���K���^���^/�����^/������0=���s����[��If�W֕�ǿ�w��v;rRh����Μ1쏫cbN��.U��$ޑ��싍�=�7�}`���>����=AUO����eS���S�L�U?�N����g�U�9�� ]�	�W�����{9�3f�6���H�8I#��Q���[� Db��]ܕ�宱g����4Hn�����>5�U�4_z�5�8�4�-Ik��2/{v��\>.|_���U}���Qf��C�����'�Zt��t7bz��[��QY������b��6OFˡ3D^#�l����#�*OTg>��6�Cw)���<tBI���i �~��V��pMAҖ:9/e�i�����P�%x�'g�A=�zN�v��+!�.')��ߵw)3�T���]�Ժ5���m�?m�7W�tm��crq}e8m�)�c�x�=�ec{�kI۴�kO���M�f	����\�f�gIf�|x0�0n"yw|[$}��ĝI���j4uR�3!����wd�w�;�sH���G?.�&3�o�OPd�d�Y�O-V.���N��������V���5��Ƨ7�''f�i�l����7�����\�-}6gU�r�=/��oG�������6g���Xw;��]��S�6�0������?�ſ���Q3�CHt_���--2��#5!�^_�F#d���d�kAwk�F��6�{qx<}����-C#�=�������GbO��\ꆘ���29�g�mM~�9/Y{�<Oa�����0����p.��C�Y-E��7�ekj�g�����*dnIk���qG3�ֻ��� ^�ɳ���q�>�ob��I �y�fu�
�hE�q��u��17[��o�[�6��i]� �s���q�t�KWe������	������v�g%#�����*���Ե����ϑ6:�7YF�Ln|�l��u��԰�{ $��3�DNc"�^npT�Q�|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*����J73��(�Qq��Y0��Ol�������O�o�=�Q�����붔�h�4�[�sF����3�}؃s�����g��<��~,�X��X����n6��j,�=�����+Q�!ߩ2q�>A�<��vl�3�Dk�{;��e�6��1�م�2�$5���=�x6���r�qϨ��p��8Z�W1��ar.X/l�Ի�=�hl�XI�I�Gn��%�M)e��_���JKF�`����s<�iY�x�U1�mMک�C�������էV�Y��ʦ&9�q9�����{�eۇsm�n�"��P�v<�Cܓr��x�����n���ߵ�;y�]��ؽ�[�R�z��z_�l��v�����,ciKJ�s���������nޝ�{V��q�f��O�%�VX�v�	�Զ�6E�U�S�gUʪ�˔j>�&��t�&��W���]O0�d�DZ^-��@�y�r\�Ri�KP�1��oӎ���n�v��iҵ���xhc���-�}�>��6j/�O�֍ET�楜�9m�Z~7�:�6�n��C%�)�m���;g�{ߚ܀�z�1�.Y���[�����`q�ڵ]O����	tq���L?}��+��G&k*��b����M���!9�Jτ��� ��qo��nܷ=/e겓n���״�V=��ٞ��Yb�fۈ�O"|`�]u��yMK��c+�2cb�����F�7W�F�5�9�^�טq��leh��:�Yֶ�4�B�z�}��wuWt�Ոm�V���6�8N��
��ũ�t���{.'M�h���}���hY2Hvi|T�x�8�b/�v^�j� Cy6K��U��?Wũ(S����R�x	s%~�n�˙]��T�6�����p�+�/P��􏬭;�%��~�~��H���s��r_�gr���q�%���Oz����3V�����g4جt��$��o���-i�ȑ�ھ��ڎ���>W�7���}�U�+B]�����������S3��&���m�v*3�'���[Ν�b6�/��i<�x�pf4�H�*a��)�=i�%�M���W�O0�o���}��9�qys{	����^{)��go�����/�A�/D���F`v�27;2)MG��KjH���i�syy��M�I�~�]���=���~�Y#�Qd�֜�˚]��9�ܞ������+5�<p���d�\��wk�-�A��d���p<�0�c� j��c�1�Ϥ�}}��&79�mZΆC lY^2x�=��6.b��N<�?E�ib�W'�k�Xo��qU�@|�U����!��6>��8w��p�}����۽7�]���w�>_��]��&�ԙ8�#�0�3�2Q�15�]L~nv򴮍�\ɛ��|��p"H���ߋ����<]���]i�l{�K�vq�/'�^I��+\���A2����nc8���m�o8���sO�ҧG���:�[N��9���:��m�a#vl9���!}�ѸZ�*���:Wc��D�ws�,�>}��I�0}����W��Q4ӌ0�i���1T�) 6^�� gi�9?R� �����r~�� �q���������K� �{;O����� �������K� �{;O����� �������K� �{;O����� ��=�7�}`��[����-�A��r<ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J����G)��j��rGC���߶ݧ�Υ���������o$�IVc<M7uoa~O'�� ��ʿ&܃_X�}i�9����]�.�N��-������Ե�U��&E�L%|�����x���˳��W��|A�Aux�ţj���ZO!��گjI0z٫&&�g�4�#kY�����ż�v�5������t�e��5�| =��C���+[֝�wzkYz�$��FѰ �,-�籒5���{�����f����U��z�-��X:���uv-ђv�ƀ�ḭ3�H����l�Q��ձ��/n��R�8X��%,s�7�ր�<�H���zf��C"�q��/�e�ԧ�f��Sv��n ��R�e��y�؝�{Z+#�bm}Uz�����*K��=��m��y�9mȟ*/H��m��{Fh�z��q��h��^��7;G�7sޒ�l��zn�f�	(d�E�T����t24wݠI���4������Q��X��L�oJ�f7������w��>%]�tu�����onř�?i���� {yv�����y�6�8����j�!�� 3C`��Z�lK��A�~��&����l�3Ij�
�vsY���`�����K��� yY���r�0>_��$�K`�����v����|}�YtO��
���{�3c����ku���xc�X��w�U���K��E�V!�\�1~��]_u>�l1���ͯh��n.Kr�����K���Z$�W��d�퍌�7.p�֟��V�7��	��7���,��]�u�������s�v<�<Դ�o'����j��#!�x�1�&�,r���Sa�%�o����R�}4ڹ>F���yQ��\d�Kj���s�^xL��	'�l�i���Z�V��^���h�8���������״y��N�Ю�maqߎ^�ɸ̄���0h��P�"ճq�Ǆr�A:)�h�-È��j��us=�l�b1@CA۔g��� 7�`�btw�n?���m,u�T��1�cNA��j�ѵ�!�;�h�mÁv��Ge���F�k��i��Ů�͸*N�[��.�T5�����:I� ���N, ���\�>���U̾��sH5,����b�������fh�8L�f�.=��z����z�`U�" """ """ """ +0�I�7�yY��M�� ���ҏ����U��ז�=\��^�(��_��]}yo���ȂR_tE�*����T���U7|}(0���vp�MXd�6���f9���P� 0�9���4��#k_Լ��p=Yؑ� ���Ō�f}�8��r����=�z�#�\ls;��8N緳����8,N���� W)���;*�jucl5kD�b���c@� %P��zD�R=DDD@D^�Qy��?wl��^o����v�*DD^!� ��ڀ��^9�;/Zw=D^n��D@DDD@DDj�/�>�������-����#�+A����~q��b���V�n;����֟�:F��k-y+��;5��d���|�����K8O�4�o��k�	3d׌������Z�c1�ct�ľ�vV�Kd`��n��F���tn��r�K��c٫X��̘0�ը�sC"��3yY��qv���Oo����i���1����`y��A;r���[E}��Y�<87��Q��<-lmᏗĴr�B�.��OLU~΁��U�-����l �r����v�ԇV�!��B\t�{�}y��C���Z\֗4�IpG!ا�G�(|Ska��R�+���q�ܒIܒI�Vg��5��?���	�<�a�'� �X�����5��?���	�<�a�'� �X�����5��?���	�<�a�'� �X�����-��?���	�<�a�'� �������-��?���	�<�a�'� �X�����5��?���	�<�a�'� �X�����5��?���Y�kjx��Q�^x�o��]��u��nݼ`�^�˚��O� ����T:�\��Rr����� �
j?"׾.�G�i|{��w<���ncܓzG������1:&ua�?m�2w\�1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ҵ��/�3�+���N�%�c0J9�'o���	�3�*##���W[���+����p���۟&�.��W/�m�qF �#-[�q?�q.$���������Դ�F��)��Q��!��l��9D��EÅܹ8p�@ߴ-¯����Ԃ��uꈇ)0�1����^F7n�.k�=���x���D��G�~j�x��W���Oƾyy����O=����kz�[$c]pj�Ԍ���s�͎��.gU�v����b�x{sߡ��I���\U�{\�l�夎`o��9H��Sa�W�_9.l�z�i�n�s(w	�ױ��߅��;��8/<��l�a��A{�R�4��
!�t��-���w��	CH��W� ��΍�\��\�q��˱W��W�l͌�YZIC�h`.;��ϑ+���7R�ZFM�0�3{So��$'�o(�-�PX��o��*�dpLn?S�k4^3rY�ut[����Oq�� ���^�e����6 ��jK���g*bbd�vc��ӏt狔�_�8��<D��b+����<�L��y�%:�ZKo��u		���a7�#�;����rh]?�(fY��q��Y�L�������,��2=���.�c�<[��.`p �A�:�G��6F���Pٷ�l<nꃷ�j� sU(��`y�M��z�G�l�D@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�}���H����ͷo�n�լ����M����+�\Z��?������.�{6������k�$���U#��.C�z]��2ڇ~�{Zl����2([�:�D��v��^��q�u���Oi�� �ZF��{J�2rr:<s�Q��A4/hk�X�0u�����o˷�ڎ��-�� �2�U:a���9�f�N8���n+��ŻO�0���gU����+�����얏Qs�qt2����f>-�[�'~·g�=�Ӄ/%���e|][h�gc������4��F����(k\[5��Q�ɑ�oW�j��L#m�K�~`��9������z1Ά���'Qdg�I�Ra���:�]d�z�.���n�`���M���î>�G;�|�la�����s������v ����kGݷ����-�W��&���vጸ=��5�4��;��^:��6�������T�p��T���E���g1[&B�\%��ւ��dr@�!]+8�xt�M|>�@ �˥�e����=E]��-9�V���6��KGo����-�!��9l�K�q�-ݨw��е�Dw߽q�cQ��f��e��/����v���9񹥤n;���XӍ���ʉ��&��Q�����f�34=�fF*��=H��՟+��|<M��f��:�|1�řk�������$�a�F�6�,:&J؞��F�q9�\��u�E&.�>���8F�����.{�c/g�qhݾ�"߉G���k������\f��ՊCH�ƽ�SL&):�+��ok �܏.z�]+��}�j'j�f;�މ�EPKjV�8x�K�y!�g?�H��oTηm��ŷ�CjM��4��nF�gm��Y�[� <�#��^��yҵ7��<�#'Ӗ��i�<��z��6.U�_Z:��9��2:V���0������<'�e�,X�&������y�m�� �Q��Ә�P�\:������t�qs�I�J�ky,��ES���Wk���8���X�o�^z���L�dƲL�3h�n*G�Ǩ�9���w�I�݇��j��o�z�`ef^94Ɋ��d"���M�ĭk�y��%����}5� �"�No���W�ӊ&2��k@ Ճ��D����f�c�d�����Æܶ?�|�Ӷ�v���iYȳL͙�LBG��[��ӟc�'��c�����/���� ��J����	9�p����Z�U4����]4�z2��W�R�fF�o��$��D@� �.w��:�������G-��
��#lq8�~D�6%�8N�ٮ�N�i$��ݤv*�TD��eU33p�/M�"�U#���l�S�_VH�DM-l�N I/k|܊�oNy�i�2����ײϯf�kk@���H+ck�/As� 9n��wKc�2���us�|aϵbi���5�E^7�m<I<���:B h�  .�-�gw��.��w\_�������2V�agtxM�~��My�s��v01��}�%�b�N���I�a�n���5�N�X鄑J[m�������=��w�Ѕ������Ih�G�j�>��z3N�s��FSe�����w��پ��H�ni�Ҙ�ni�҈�o\�u�,����x&c ��;v�=������ �F�df�y�]*QӸ�����Ļ%;�\K+�����I�	��ٲ�`�f��#�C�ʮ���m�k������Ò����b0�~�.��1��fj���iUǶ)�,ll<V6wYË�9�l��,��� Q_���jX��z���!�l�����5�pK@ ;nC�鍩%t���W{g��Ϥ�������qJ���ZĐv�rcsI��Eץ���&���_b�U��L{<�e���$l����~�����;.�n��5v>&M#��d.v�oW�C�<^�c��y^L����V�r^��wDϙ��;r��e��t�%�Fd�s��y��Y���ؽ^��""5|�YZw�K����W�~�����}��8��1姇��c>K�
+X����>5>�3��!�������݁�yT������,_P.	�yt�Ky�OI�V+����ul�g�{��=�dk�ߞ]�2������Ә�y�n�:U!�ŉ���E��ǻ�&�������Ū��S��K��a�C5o@�*��l��t6�Yy�x�af��8�ҷ�}K�k��>/#������a��ڷܯ��,1��$Bw<w��G�!ۼj"���\���N��1R�������:F���A�!�.Y[��ڿ5��7�Ķ�,���Y�H%�ВZd3�x]���k:cU��Xn�����j��'��\�هg�xu`csg�ܘ�g`9���l&���I�C��׽->����]dm�=�3�1
[��Ěg�1�+�j�M_[5'�\d��u����e�`���7g���6�V�t���oNM^η���˓���ܯ�$|B�]S^�� �x9n���A��g;GOc�{%j*T��1�L��=�����!gq/����1�zB�޳�����1�^�Do�=��;v�6P�=����V*��KZ�_�^oQ�쵙V�Z�2i����=҈K�8Hk y�	ߚ��'���g1�s6C'r4��<�kG��ɾū���ʷQ��2Xr:�3��b>���6��gp�y<�ؑ�־��>���4�[O��uq7M�u�[��oW#�����o�]{Q~�6�q�.��صU�c8w-�p:֬��r���F���p�8�
y|��\�}Yӥ��:�f���n:\��22�ĵ�Nܻ���}J
���X��� 
io��{�F""�v�����<�e�3��>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��T�j�=�K�-y�г�7uoax�=�IO��Z�olf�wa����&�q6>�Q���q9�����\e�r�j[V�,��i�`��vo�w3����m�}���δ�-��9�Y*г���]<S��k�� Z6 9�Ͱ�ߗD��X� � ��#�pe�d3�4��cl"`$���w'�<�Ku�#e"t�M7�1���r�ԁ�Iz�����;��I���¤rN%"�T�h9 �;�s^ﲌ�Qy���E#�E��=D^ �y�Q�|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*����K��!���>7G�6�a���F�GN���g�!�� t?ti�c���w��9���zܹ�~Ǫ6��19L��+cێ�z���������Q���m�2�~8of�/�3��捕鮪?�ZQr�?�_?k·r4�X\v&�l�ۓݻg^8&{�"0�ҳv9�pq�߼`ش���^��ݳ�2��Lu�m.�lmJ�Q=���.�a˗�W�V��L�Z�d�ա�Ҩ8-pp�޽��＀�n9���S`Ƭ�D�9oy �b��9*p=� �!�!��<G�]1]U��}]1]u�3��t�FU�����I1��c��0�K,R�1��n��/fZX�� g[40>F3������CR��L���J�A� %-q.{	p#��!�;.:�����j���}u�в���ۆ���=l\7�k+6I&������o�xX;�B����S1Ү��3�� ���3CM����㛿��w��ż��*��q'�����3���sR�'���2��;�Q����D��p<�w>cŲ��Zj�.�Ϝm�`��񴮶���2I<���q�����{���ʥ�IbZ��
���!�NIe���FX��y8��<�>b�Ubr*E�o�xN��¤^o��Y��H���s��r_�g�􏬭;�%��~�6�=���[�'�h� �x љi� �k?@��o�+O����V���-��_�9a��2�[2������g0�}�݃ym�(7A�o��V?�{2�}�g���wU��t����(�RٌK~I���/�1��۝�q`#���j�g���w��u�|qڮ�����ݱC wa�.v��v�s�(:�̳�V��� �^{0��V��� �\�ӳuG�SOZ�"8��_VD���Fozw�F��W������~_\u<Q��Al�3���A�0I#c��}�b���?����מ̰���g���W��+kKfY���U�V�]��O+��&EH�#$@��F�7k�<��k+�c��!�{�c�v�$��g�W� �{0��l��� 5!���y�n�����׎�1��հG��� ���yl<�[2q�6e;F�����o�W� ���yl<���-�V��� �Of[����� �6@� D���o�W� �{2��l��� 5!���y� f[����� �9��-g�����-c'�lbn�J\M��<� ��㉖F�7�dm���7�A=N�w�C���f<lB乏rM�X.�L���t�9�f������ �7��\�1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ҡ�YY��q��v���L&^>�����o�_���?ңo׫b�<�(d��e���;�{O/z� ���)3/C+b���ųĜ!�hq� v�oڷ*���R��U�ۚN�e��\��`i%�;x�'~|��U�4_z�T\�@��S3z��ll�)�<��ղَѹ�qsKvk�{H���ȷ�7�u�P�Oc23ޫ^�6d�h��ܛ�-������sC�͹�֔M1��M1�惎����	��S��.Y���C����`��� o�^�@�;�55��ޖ�+�����"{�q�V��ԶVǷ|�w=��;nVŋ�Na���0ױ5l}�z�-[�~�b״���'����;��a��!�qE�V�F���8�2D���4�r��޳���OX�Η��(�[0���Eb�,R��ϊ�&H_�r��jT�G���L�_V*O�N��e����A�൥��ͤrX�^�E}O�3�a��VS�n���8�[�%�������)�/���B+m����K�O=�X�W��缗���:��F)�ι��GW>铦{�g���mLu�,Vt�֝i2�(� i�s���Ҥ1��R��k�9�,�଻���*��O�&"NN����+u�i^f�v����gU��� :�D��ܞֻ����	�n��u�=�����d�(\[�]EŌ$r%��[�lp��x���r�V����Ai񒒴�e��j5��C]5��d13sɠ�A�=�sϱkZ�P�J�|�p��V�{���K/i���vw�����ݵ&����<ؼ�fڥ)c�	--sǵ���5�k��P^��9�V/rlĵ���ͱ'Z���8��{��ĸ�kz[�{�Zպ6c�֪�kF8c)u)\��y3N�3�v����\��/5���{<�S�n�vݾEG��eH�#%��hJ���+�����cK{��+c1�۱��_:�E�m�2�d���c�g/�\-�+VuCjfێ~3$��ֲ�u��s���;��ܗ <@��N� 6�o�A���m{��5��h̓�ێA�ˉ�y@s�%��kAۉ�\[�8�;������=Ѷo?�3�%���,� ��0��K������n�F/��d��m�|7���*�'�(��^��a%Ēc'r�b�"��=[)�j����n[]X�3ۼ�q�,$p�ό���'�|���Z�Q9�����Q������$n<��fv-z����Wb�F�qe�8N�C/U�$��^�6"I;u���QY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�AbvւI^ZƗƗ��d����x�Vԕ�a���>��v.~�m��7>e��Ϧ/~:�`�j�.�9�qlǋvﳇ y��; �q�{3��v3�� T~3qf}�x�ޗ)恓�$���ׂ6�6h�ñ]'eo�qm��!�5x:Q�6�{2/5��{�[uY�]��xlŜ!���w�+xu�m�N�>ȋ����U%�,/���c�{�x| #m�B�����2�r\ݙ�����1�Ts��wl�n�A�.�՗�4�J܈�6[���G�;�>���j��~�7����HG�N���U����,U��mI��>8\��p�=񽣈�ad鞐���Vg�t�܊�.a�ˏ�8�<y�G04�q�=�h�sZ�#�f{2�'�ci>i�>s�3�v�Ґ}�ߊ�o�j��^��l��c�v���<?�{V�g�H���ifc�R��z͗h�$���G�As�݃s�c�3:{��^��Z���8�6ԇb�q�w�o�� `-�?���9j0dj8��F7�o�G��aE� ��=a���lY9��29�5��X��v��PLMz�y�1�y������δ�/ҷ�F5��#��Vm�ׂf��F^�À�&�͹q7��o-�R�U�{<n��a��8lH>#�kz'@�F�Ԇ���4P��TȚpozѱw|wq�vDc^��c�7�Ε�ts��)�d���X�Î{���˶{�������UK���q�,t���dY �}��gs;xxZ����6�&��z'���M9;�d�3a�������q�'lG�*�^�k���eBwԆ��qPs[��N���8��n<��n�T��.� .�����u���^c�q��< H@n9�cq�Y�Lř��Û���:��WmPxY[�p�@��Xaw�"@���v�oQ��􏬭;�%��~�~��H���s��r_�gh��!��e��d���09������B�p�{Pp�H�����`�*�L�,���vq^&4�9��` $���+#�,� ����o�A�[M�s�
��`͋Pp�H��]��@v���;�y�M���ˆ�bF�#L����	��w�;�ە�b��3Ūs	�$�� �A�#�V_�Ԣ�xX`�z|�$$�8Gy����s�?"dk౵䫳��=������f�:�YdlQ1��{��h�$�o���� X��d�~>�xK�߅ނyx�(5�i��S��L�4Hݤ�w� ��qnAn���"١�$�8�H�0�������!�M�N��~��wl� �����V^�ʛ���?�2�&� ��� ��7���ي�2M4��(�s�{�Z�;I'�*�#^�Z��y�<h1;�ĥ�M�+���~����(ܦ��alAC'N�ӝ����c���S3���:�� v����I��;��e�M�+,8��f'v����I��;��e�M�+1a�l� �����U&����_��ⳑVK%�O$}P�kI����9�rM�X.ȸ�cܓzG�:�3�mO�3�T��;�U8Ͻ�?4�PUS�?��YA�?��@�F�cn(�״�,����V��8��^u=?��A��f1Fb�Ks����U#�}��>t�+�ľ�V�3k�D��=�L^�^͹�A�e����/�=KO���͔�E<�ا]��Hظ	��\;O ���>e�U�4_z�]T�^���Y^�m����71~� �p��� ����9l{U������5tt͗����zS����۱-��º1<1\7��c��ږ��7�mI�u;]i�F3J���i�\tOo`< F��߷�g.�nKp�o[yW����i5mU�i]du����r)_a�[��݀�����`.ajW:V�j^�uݺ@�3zz��	+��\ �A�0 �Ao�c�TŪ�1j�v-�t;�c�J�����8���c:]���������C��J�$q�@%�1�n���;���M���<�M���S���{��q�w��7*�����t<r��fQ���FXHt���`�HP�O/�Һg36��d����XXθ�״� ב�.�	�^l�ai�\u�U	��s���3uc��9����6��4��}��7~-��m�t0F�9�i�ʪf���y��UQy�Qy�o�QY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�Abb	#.{�L;8z�s��$�J�I�?w���q���l�ѷ�f���]�¼JZ����}ơl��}\%\���Ca����:�I۳Ğ|�A�b�<���q� ��@����{���g��<����6�C�=��,t*ܖQk')�6�o	��h�;�#�;	
6�z��� @[�K����a�e�V@A���4������?�v����<�n�0E�cn��9-b��q��r"�a�H������u���*�X�Z�#uh6���<-��K^]�	!n=j�vl���!������{8ZHy��`pqp�; ߞ�6�t��e��iYC׺��T������I���٤�Wq=#���kA<�Y�q�[VzϊV��L�c�-=X.��o*��S1�����N"�.�����U��&��6a��*L���p<8� I���n�����tɬ�7��0a����l|A�,x`p}���ܩH�jѶ�E.�,�*әEIK"�į�=�;09�s�R�o�*Z�Ug���ނ�&f�,�U{"��l'�c�����J7��W��q��7�c��}w���k�$ö(�����m��w�v��>�?��#����.����c�ӽ���<d40��a�κ^��Xm9��sV�Z��v2nfg��ky���{�	�V5U&AK|nI�����c�<܁Ű<=��v;{,1�,��Ft���t�q���c%B�%���	U7o2ַrK]��n�����i�'�}�cD��U���/p�|��M��A�r����\D
�:WC��-H���$֭�w5��/���[�v�L�Y�t�*|�#�uY�fM6X�s� ��Z[����|��Ë�zJպgLg�K&��^L�O#�_lWB�����kb;G��u۴����!���Sϊ����nLi&�^b	_nRN��"6��q?~кŮ��m,g->G����Ϙ�]Z@���t����<A�tRݸ�ogbɩ�Ɨ��n"r:��ˏi5d��!2������v�� ���1�j<�V|V��;%�9�˙�v�M9��D��;�մ�"\7�J�tU����sX�����b9�ָ��>���ѧH�Ηp9+uq�*ׯ~�.H�Ws����8�@�Ûw��SZ�X��Lx�e/��6ԭ�%����7 �ލ��ŸU�<��;{
��3�8=��sN��@i}X�Ek=��c݋�i�3��(� ��$�^}����'�.6�y*PZ�H"�����v���lA������������������_�G�V���Ò��?tſU�_�}eh9�|9/�3�LA�9ˠ�� �����ش��W[M鼁�����#t.�{]	iih �D�^E�uͳ��� ��� ���}+Y��U�B����ݭ�!t�{��1���ej�f�A�ESNbj�.Jͧ��3g�du�����s��̜��ݛr;��M�Ka��Ⱦ݉,K4-g;��H�`6<�-�s!���S����h3�wtc�����X�s�K!�߮�n�gv�bfں|��n:�b�\q��)�'Cج�%��[� �TG���驜�"t�{c����q� ;I>%o����3G�s�]���z]��yyx�(9oD2�5v/[VW��9YRT��#�����=d��� ����(�n+��%�=4�oU�$���1�٬�dL/t`9�l؏���s�6�6n�-(��3�5�e�S8M�e�۾3^H��q7���%����5�]���~;)��{uod��d�Zv�aa���S��Aiis]�����6/CynP|�h�̦�u�+�l^�����\�al�Vw�������w
RL޶���=��#�f�Bz���aZZ�e�8��.<<�t� �{����5�b��KVd3��RP���ޫS��31\�$veuο`X�G���9r;lW��gI=&}����=��&ls������ -�f����_c`t�#K�4x�|3���[�a���"�tL{�s�;	�4���U5Dg.-V����h���x��4�mC�{+P$l�y7%�v�0��ˠ��6�h>�V�p�k:f��ﺐi�.{�Mu�s�7E�b�"��㒤DY�q�ǹ&�d\o1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ң���w��1�d��<p9��x��;��B� J���k-���iΖA���+~n'7��U	(��Fhd-{�+b�<����'n{�������Թ���d1W��r��a�؁{�F��;�>�g�����I��h� � ���Z��i��[�Ԗi�.u�e{e�CxK� q;m�-�ݫm^�&c�bf:4�1ZC�r��O���#��>ÃxX�����<�����]1SO���6;��Zn�V��9��o�ݮ�ۘW:X�vu�����i���H����i�i���V���'�f��	��rY��cū򹎭4rH�J�w2�������ޫ�;�z�k�髹��P�����D��trǳ��X]ð�w-�nV8��I?���oO%�v��$�fp ��q��b{�s]jl�S���=��3�ɋ��$���k89p���;��.Ņ�,��յ,�B��7/�����]����Hh�����ݻ �w��N�]2�-E�����]<����F�o3K+�!Nw`do;������7NǪ-Y���q7$����ǎ���o���k\gEvl3��v6_��ٷl?��J��ȣݽ�c�����@
j^�J7sQci�\���[h���=�,���A����ʱUQ�QLs�kw:>�kf���\%ax6XrG��ZR�h�09����ۅ��#���WI��<�����f�3,�ƶGI�ư��A�Nq o�j����FcD�q2
ػO�?'QhL٣u�Lb[Dmp$vm�Ji�{K���f�w-�O���}wż,`�iw 6;J�]�)�W��1��L�5��`���r<�s��]��.��m���w���+a�T��ˆd��"��/ۛC\��7����]���e��dE~H���xKA߷�q���t=�iu�*���Ё�.� ]�����Hz���<}���iM4��\�UV}]��
��4l<�9�vv�oWt��My�hx��߳иu��s��9S)9�ߖ���1��NNK������n�v�ҝ�߫2ԍJ�:�G+���X�z��<4�N�l�nb����g����4�Hό�+r\�&�Ϛ65�g8 ��>Nլ�?��8C������a��Y��D�ƹ�8�s%��l��!iN��;.'!O��?!6K+��Å[|}[^Xw����7��]�4�L�fW��'�:^sTc��8�ۜ5�IL ��G���x��Ռf��fr�1��	�Wl����Z!������G%εF��n;cq��Oc^��9�w<�|��;��9[��l���4g��5b�w�q� q�N知MQE4�'2���y�V�V�M�����ḓ}�����+$Jл��7F夛
�v�|��{>�$� ��m���ܭ�M�XD�9�V�������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J#صK�;���M٢��m�#�ؼ8����ff��9�c^����Zῐ�`�m�G���J�>H"��	�#��q���Ű�o�(:F-�6'������H��$�)-�=\}��)��='e`ً���������]�3�T�m>0�`�jԳ$��D�:�փwtR Iܖ� gm�!G���g3ܑ�)�3Gy�����ֵ�o�]���m�b*o�i�O���X�YL������N9�-�9���Q�3�����@
Ӻ��mѨ2-��$2�ˈ��/s�6Ŝ=Q�ۇ�ڵo��YNMrʶd�_��Ў(X+E��6=�a����	#ȷ�������P�,�YZx��G����أoqp��ͼ{�V���U���y�����|=�{29	�n�:���/�4�F��{\�\�m�ߌ���2��2V:���ǹ���ֱ�p���6��̶4X�Gf��;Q��G)J�G�L6#n��|cʢ��Ν����[!-6�A=�	�cA� ���G���Q-�|Y*i�h|"t27����Z,}��x��&J�q��cfFB%��Z�#��-<aۂWDDcU}�X�S�sX�j�1��^�f,�a2]����	⌆���b�c�{Cl\�d�j	�cv�餫5b�w��6w��{-�jz��z?�+V��61�2�Q԰Eilؖ��-t�<��v �rXJY�\]��畳G��^;Y肀�Ѱy�����"l媒9�rs�Q���,����0|}�L��K�*+��G��/��c��؎�M�1��D�I/�s[������,""" """ """ ""5|�YZw�K����W�~�����}��8��1~í�C�a� �W-�f�������	�q9��
�H��z���;�`��ݖ7��&�?���A�u;w��R�%�nSu�CN��qcy7���s+\�կc↖�l8j����i�{OM��I�����\I0{�6ۑ]KF� ��\�S7b,t�Z�l��"(���q� ���[Rbu4�����7p=�e5��}�=�p�S�u�Zܸ����{���;�"Ls߻!���~��}���Q�k:�|��e�L�,TQK�:.���8��%�����ws�ۊM�=���B�*�����W��K&�𱠗�3�%��M��� �7���
=����l9r���{vyy �Z-��Gڸ�Y3�8�2\$t�s�Ǝ("�qp��1�V��d:;��N,�W$�i�X� ;þH�/!���0�O0�_J޿[J{�'��Hd�y�����'��X׵+f�{y�g���9fk].�k'��{6�5����cD?$̛E�4���4���.:Bb�#m�ѹ�;���Z�Eڋ����7)͏�bq����5�5A�:6�-l�M��Fm�>_���U�f�xlG,�\�O�qhp���y��+�d��GtE�q�}_���������o"M���o�	�-^vC#�l�\�A����̷Zk���Z���o�n���!W)��#���$�|2�1^H�RJ�E+�ps"v�Ob�:�Wa�F%�,�����Cz�?����7� �����^ֳ6 ˂��)��s$���.c�p=��į�Tӽ�L��ong�����ä31U�f���)ӻܱ=�j{7^�4v't$�?s��}��!�4FK���ye�6�����k�.r��]<7p�*��Y��5s�/�S�E~�e�����0���\;>E���̃��6�bw�#�����W��X�?��5tr^��W:����a�itq�����������""�y�rM�X.ȸ�cܓzG�:�3�mO�3�T��;�U8Ͻ�?4�PUS�?��YA�?��Ae�\���G��;S�	Y���dx �� �r�Ƨg����˶1��H�Km1�d��;���p=#��k�SQ��d-Ӿ�U�����s�c��z6w���}����c�1��u	 �w�1�����~~���������Ԃ���/W����o5��T�0olV�+�l�=��ܱ���vr�n��[ҽ�����gv���'�Bcl��8���Hq�BF�`9nN�r�6ޚ��f~����fF�@�L�{�A� �����
�%��:�*�^�M�5�l��'��v���v���>�c�ckZ�J���P��  �t�~�u�.>ӷ;�f�s4�1�̏(gd���'n�l./�� :���܇4��[5��,�f�=O��fN'�c����� �۞��v��zb�0\2��{&)�D�G��6w�9�n�t��2��d�ԖXa��g����A�ṛ;na����?W�+�J7�<��-�;�Y(��X��a��=�'���d_��h?NP�:�C/[��)ر�iq-��~=�N�:=3���]q��{/�l��ËxK�w�H�N��B��/sB�H4��f�JfIdk��h���x�����f?Yɛ���W��6NY������u�8���v��Z$�9)G.��:b�Fֺ(f�D��[ͧq��_����~��`�ǰ�̮�@������O}����#�U���(ꌗ\�Y�HC�Csm�� ������߉ý�nOj����\�Ơ���I*Z�����U�óDfN�G�l�K���/�"�ᙨ��ziYc+,�-]���nk6ld�ƴ5�r=��rw7�gэ��w���5�4���b�T�.ҹs�2p�
�V��n|]on��|{��X�1���u�o���|Ek��:X���]���Վ ��cx�.��:���mY^���S�yȤ�n�;�s7o�aoa��:
�؝E���m���>�dcjEfAN�qoK�v'�a�h׺��KY�>�C^�pi�i�d17��h/����7>%�4�L:�|���[�׹����Lq�V�Z}dq���7`'���V�fv[r��Ʋ���cj[�yq��lv#����in���b��)עr_xx�7Vȝ#�v����\�Ű�S3�!�j���J���ONX�B�V���D|z�KT<p��=��݌d��a�hn����-`[��������=��T�l�h`v������%��9�-F��U���Pt@T��2Spo{8� ��N�n�������i��X��*Y�e�sb�j��͒`+^�����=��)�1����ft��_����W2�|�G��uY'�"|�Dӓ$�.�h���p�w �k:����J{��c��c�d��C~�gH�!^�Լ��9���$�6
Zv���j����6ܯ^'�x;�`�2�v�nݪb�F�f��f���Ĵ�(�+�Ic�ƿs߆�r�ؒTc�Vj�����a�^8���˼@� ;�A�iv�����kS�ɨ��MC5]=N�{6=��6D�Ei�k]�"�8nAo÷r���m���Y��hɑ��:ƙ	!��fo�C����o57�l�������lUoL����I�rۘLJ2�5�NV�G���f�f&�r�㤞�� ���X�w�8F9{`���H9=S�u&�
8q8K��c#5�%{�N������ma�;�mÿ=��M5�����i���V�'ypi ��n�ؒ�� �xƻ5"�x��R^�f�V�����z�ׇC"���Gz��GN�/��D:�Sa*׻��b�݊+R���8����v�m��~��jյ�J:�Gf�>��V����,|9�&C37|rA����ւI�`N�����:�WY�Xk��Rz�z���x����a;�F��ϱ\=h��
g�+�kW��a��t�rs�|e�G���n�H;�)_ge�[ZD�2p9�n6|okC����-�}��l[�ڍ�s�u�l`yI#��go5���k#��t9#g!M�Qe^�Y�ލ��]� ����+���et�2X���
�7�&]jP�c��X@���pho��Mک��OFܽXl�j�K`<�I���#~��o�nB���|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*������{���#i ��9�fMuUqrIU%ֺG5�X��pi�����{�gEך�j�b&��qg�F㻘��ٸ��΃g��l�۳���,򣱀G<�`�?�RCʠx�9��}�^���u���U��^�b+t���a���#7k�G" ���AҮz9\��bq�C&M����<����� G!�n[����p�+U*7�j^�y����X�lr׷�;�� |{�*����X�9�,����9}��2u]]'>N��'�	7���<Ac��8�'�*5���������9��gU�p�'�`�?o4B�;�[6�2ܐu5lK3j���;2�(�x��Ǜn|����
=I���Fbr5]��B�sŴ28���;�6�k^����\6"�:,�FX�R��|���?���M����t�'��kk��Ê�9\�[m�&��،V���pu����|{n�/S��N�����T�i[^����v�1���{�ǐ�'ı��ve7;��C�{�o���r>=��J尔sԟO%N�_���>}��n���:��VѪ�$��3�$ �ny˟$6l�R��� ��^����7$� rӡ�s.��[')��}e75��/�����|\�'`�z�Y*V*X`���)������ �l�MÇ�T�����Y����c���Ȉ���և�	˝:�:�bŻU�bl�r,uw	+�]�6`[���C ��r�Bʧ�������������+���>�p�wBמE�[�� {�Z���0��Nd��9�M��n��k��#�=��!��G�Ն���䶦t?���*طo��g��Q�&l��5b�w��6w��p9��ފ�P��L5�lU�\UrWq�]f�GV�5g9�ǻ�$��s[�{Z�)Z�����ۗ�G#n|m셜�tl�*Kby,O����,�v�s��a�䦲�s�rT+�l.�X�?��Q����ߗ����T���~	h>��W�=� {�Tr�;7vs���6 6y5=>�L��5%q����]��Z�,����6�iE'9�$1����^�#�&L����X���sO0|�-Gi���aq�e-��F8�6���,��9����vR(���������������,��_�}eh9�|9/�3�L[�_�G�V���Ò��?t����?A� �W-��U����2hlF���$3ן�{W�H#�	ީ:E���7� �����[�?IX|TF|��-�^&��/ycv �����EdtNoYؤo��IZ��?�rT�GO# lڮ� ��y��Ⱥ�0T�z�fps�#�4��{�ܹĞeg�L� ���;�����эx��0Ks�ZD���q~����;rwX���[[#���9�r�8"����e,��m�d�6q���Y�	���?tM����N��#��A̺З�x<�<�{+�G�l�f9[+��nO78��-U�����f��2�M�]l\r��ό��d��ǐ�Q��Oik7<�ߺ'�Q�H �0� �G}0��\��9�u�S9�ľ�?"�R������A	�1�%����pozw߲��l�����1�!z�J��L�X�#�6^	>)�'ngm�+�wD� �;��tN���L �?d�F��w��W0��ӱfz����Fvܵ�!�#n�ۺ���.����ƭ�V�'����lr��񸹌s�CN�o>`��޺��w�ξr=��lk.E�����:;s���gb�b3��W}0��� w�����V/t��U�L't�����A�����U�L/{��]���X��?��a;����aR�y�rM�X.�l�����\�.w�7�}`��c>����=AUO����eS���S�L�U?�N����g�V���=��X�:Ii��&��s]�wp!��;o�`[<���m��0W���\@��O��;�p{�/�v�ܟI�5�V��R���;аr��|��x�J�ח�#��vm�}���S3�8��wM��d��	��{��lW�M?����������	�n7#Ⱥ^��l�zc%��'N�P:cN����[�Un�g��y�zX�6������ʏ����7�A�ii�'�Z~C������=��)�<Tm�nwZ�Y��w#��wܞ[��w��$���Lm�}y�62PҧP]� W�zn������1ܸw��9�W}���6�б�|���G��?���7�?��=��b�\��R���5�28܆>9h��vNvd���6����Q�޲33y��̀[���#�ޮ"�>J��0թVY�,��)��v�nͶ��Q�zc��rx���M���e�8xem���uGNKx�p��۸<��]�t~_�����l}X�����R��ݼ�)���J�TLe�ҹl��;(�f6k��=�i�`�p>2��'W̃�v-���V�йH��v�ے~G��{��t\�[÷߷����[n��?Qi�y)`5�;K�E����#�V1��M�6c��C���._%R���U$�>'��Cf�ۊ79��%�s�5^�U\��UqLf[�+BɄ�$0�̌T��c �3ٱ#��H;��ѫ��	,�c�oY<`���c�aZwE��!�૏��e|�������6h���o��v��6%Nkl��d8wU��f�V�M���?g7���h�k�s[��-?�J��:��4���d�X݆�m�N�����}j<�KJ�7J�GP��B�.:V����9�K@?q'���m��v[���+�-cK����n�:K��#��*�ufc�e���g��g[�m74�����[QU~JU���}jl~��T�=9��U5!;[��+���	;��d#�܇�`����Ɯ>@��5k��/q�h�l8�.ݹ�?ғ�ɷo�֘.��e�(���"x\Z8����m�%	����R1o�ōm�Uy������d�3��k�h<�.cȯT]���V&�z7M1�Y�o�i���Y��Z�@nA�x�a�x��3�->��ׯQ��b79�Ն=�4���;<0;� ����G��;��j�jS��� 5�9�١��,o�����!ki�E:s�A׌��Rp�7��JG� <�(���1�~SKIgGz�ŭ�2�7#-IoZ9��+Xt����䳁���p�=�ߣ���5�������v+�I����4���;i<\|��[.&��L+�P�K�7V�p��m�ָm�c��� �\1�֦��}cG)�����&���At�8�7��gW n���f'-��{1
~���,Yљ(�����f0O~�[F����Rj]QW�e\.wr�fs��d��k�	-o2�F�r#�V偎�|.><��ϓmx�fX�$�4q��'r�&�ݖ�9��=9��q4uGtT�=̵볉��=��ݼ�n�:�*ta��Ѿgzds>xf��2��`��pl��]�f�E��y�x��ZI���}Cl����h��<<G�7�uƴ�Iz���:�ry�~fJ���#���hk�i� ��x��.��8J����[�hF�>ey,�?�l��o�=O�t_z�g��������f̛�����Yc#=��A��KO!�N䀷栽��i(g�Ɯ��U��읣ws� �g~߹�����Z�=6�Om�0�V:���fY㐈����&����8v�Qc���:�5)��a�C��28�#o4�s���A��1Qm�Zleǭ|q�N�kZ���j�t��~�Mv�9�ׂ�'�[�����6n��nxw9��� [� �����ur��G9��B�`m%S<a����|�=�7�g��vFx�8:�B��t48ᒯ��iakb��l�{mI7L��ݏ�g���[>'X�z�7������D�b���{��Y(��0���;�y�Z��b�_���j���
��G��bA&�;���O	!ї��G �&�UF�DN[λ�I�t�q�G7#Q�1���$� [#w'Ȣ4�ܖKOҵ��^��bk�ʳY�o�qc{|�r�^�����x���145m6����G�=h&c���wp�'��<��9�ԗ��<;q�$v�"�+0�I�7�yY��M�� ���ҏ����U��ז�=\��^�(��_��]}yo���ȂR_tE�*����T���U7|}(#�@�U��{[#KIc�]��G1�H8v^�8ZSR|��wR&���É{�<�z݁򐷋|pH���^-�}����-k�SB��1�����8o6�Ɲ���]�6� �i�ym �ܾ~��K���yFd�uf؆Lݤ6��$�G�浢.�p�H���&7��9>63���y-h���j.nD�'#��x�͌t�j	��l��L�-H��a�]�o)w���;����CwOt9�1y�~��y�'G#ac\���}�O��MT��5]���¡ؽ^��ŀ���" """ ""6^p����􏬭;�%��~�~��H���s��r_�gqӇ� w�%��"O5��k�d=T��U٘j�#`��&�����l|���wAY~��|���Wf۹iE	d������ZŬۛ��_.y�v-by�:OP��΍��J.��fv�]�nۑ�j����t��կF���V���! �;�=5���O�o]�շv�:WV�4-t��9�7��ȴ�E&#_�/W�T��qf䖕h�nNK���6-h`'n}�浢�5ѽ��sSU����Cn���P������O�W���X;�c�	#�v?2��I��\c����t��f�dFؘEɞג�ǿ܇V9t���u�r�cTg����goi�3�l���:G��4���;�܅x���2�u���>��v��V��d��n1��l����[���棹������ۻohD�r���ѵ�s	c�p��ȁ�\+E�ژN��j��$���XnJ�otY�y�o�˻[�6sZy��
�i���=�YME^U~���_����ڞ*�7�K3�Z=$�!�R�8$��2��2@D�b{ӿ>@�y+��[R[�5��wd�[�k�L�lg�7����7ߟ�h�c#�����x��$���As���7q��߷z����v��X����4��p�n�r}/��7/�tnYg���O�.jzV_h�"�8�c�y��}�k3�N��s?� ���kۥ��kX��8c|�4nv�-Q����#]D�� c���tY�f-֣�l6�~cb��Yr�x�$�ll˜v���c^^��#T��\7���;��g�� �-���=i��gBt���e���"�N7�	��:F��������#IT�FYNЦ"y~�x�'%�՚���e^��v:=!���h�s�29�yt��m�6f�ʻ��z�Rg��Pg�.�V�|m�����Q&G���.��ϒ˻Ռ�ki��9���'\���Q��f2���Vݫ���`ӽ}d|\@���x_��6m�\�L�=E�u��c7�e�W㭺(k������$s߰<d���hk�UT�� ?Unk�ۢ���Y�k��Z7B:�!�z,���ϐ�_y[��Ů-������r�WtM����F�qr��<�����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�x� h�AXٌQC����V���Z�ϱwn�-����#�dI���+V�c;��i\�m��ň��~WDǲh�K����Z�÷1��v�L�8&2��h�GPAr��yb*�V7ǴQ��u �p��g"�4�������Lik���W�!�����Z�|��_?�k�F��ըiIc�#�Q�����$d�X���w9-�@�g2�2O�.ˬ/X�K�4�|Fk>N���z�P�b%�b�Nǳ�զ��yʱLC/F�
9ڵ��G��bj㤌V|��9��lHi��pG0���h����xc�Lg�qb6m�n�@<���s���A��>�ng5Q�8���&k(>�l�u^���� ��5�^�u,,��̵O6L�a�ۑ�Ce��S��`���A�&�^��z;~"!b�c���K6/�ic{�GH�� Ü�$>W8�\KC�wG�����B#GU�s6�	!�պ�������q��o�]WL�29Ll�2x� c,wL�xq�+����5�x��U��T���w�d.�djc�+�qS6 ��Ʒ��ϙA�1;%���bg�F�Y�)��3X��繤��C���G�D��!���1z�G��O�%<�ΈB+f��7���b݆��l���Cyl���1�6�F�K�F9���k:�,�ہ�[�q� 8|jbf:���8��SE�#�f&)#��sdd`��Fw'��v�.Go�ֺ�J�y�-M����OJW�g�G�&�v�m�ϳ��e��~����j�[_V	d�H�%���o�iۑ{T�z"�b���⭌�k�r�)ؕ�B�,:����X@�ɤnݼ陙̘����stR2�:>�� ��� ���*���4��'^�:����w!��1�p����-���
ʽRk��#b-��$��ȗ7�0ԟ@T�7�;2�O�f�����Zkcl;aȼ0燇s����&!jn����K��%Z�s��6k���������z�&�p:H%tm� _R��ٷ��y��t�ί�W���Zw����V�nlM��F�yN�sRdn�/Us>f!K�f�]����>w��R����e/�#^\�yA2I���+c(�&c�����6��i�e�Jq���Av�v�n|�`�k-�`���	�?+�&?��{�t{�x�;y�����33�=���F�Hֹ�9�n�(��7Kc2�x��Ij�0�=��$y��T� ����y�쳋�f��^0ORv#v�ď�*�}��A�Y��3r�{r����],���yT� ��1P�2��}q��#��J]���4��Gۖ�_����J�-��M�0N�5�����0��jұnx+G�$�# W���)�h�^+@��#/��"�v�o��\�}���vs+aDt�KJ�j�w=wJ��ah�����$�˾���.D2���Lmj����'jK��g�b�$��k��ַ�6(� LdDx=+_��ߊi籘��s���ka��������Ǵ��Df	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�Z��V�Z����ȣt'��w��q��ۘ�]�z���8�5�-<.-;!��Eߵ�8������1J��`�@@;�H������bp;��!���Bi�=� V�ϟ�\�:P��e�LdkG,u�$`���2I���X6cX<��Z(މ��6�n+���>�.~|�&'/O=����؎�Q6x,D��$n�����rX=_K;j�����!�Jan��|n�\�z��#g6A���-P����U���K��)A%H������,�#������m)���h��4�y�݋�N����vK-W��cN�7� |���� z���@�;����/�e�_f�ts[2�b5Aqn��͛�Ti�V�ӹ�9J����K�IZ��m��8����K��N$��AS��x1�v��}l�\T��B�n���=���z7
@�0�l0�z;�-��Y�V���@��|�5����F��ߖʎ�����.��9K���5�/uiat���y���l|�6�l	'��c�&�c9v��^�6�X9�D@DDD@DDD@DDD@DDD@DDD@DDj�/�>�������-����#�+A����~q��b�N����|�/����F`������#�X�s��w�d�/G�~�Q�NgKPc,�5�n���A�^��
���u��D4���^e6�@&f�[{6nC���^��p�0��^����h�c��4SWXB�5����9L+��pu��������خ��Z{#%�Y�ՙ�`���8�FûG����)of(�7�	����a[~�UxTzCNi,>����||8��#�v�w��O�BO�抱����n��$�c0�gu��\Cnø�p��e��7�	����aDWTNbI�D�D�F��X}]DS���k5�Md���>Q�>p�q�i�L4"���Z:2�z͍�ur9��p�H�L{/G�~�Oe��7�	U��m�3��h�:#��$T�A�,|tx�s��g�7
>�D�B�>���)*T�I����#{���<�D�|�b�b��p�0����n�~���tLbaW�}3J(�R8���-`��<����$��X�ފ4�"��������e�����Hk���[�����b��p�0�~�Tp��o�M}�cNјP�E[��~���� ���f���c);q�	2�kn��~�5�=��г}����?L'�����z�-�H�3�p8O�..�8ϷXan��v|�s�kZ��]�s6ry+_j�i�"���i�cC_� �%��/G�~�Oe��7�
�ݹL暹�U�uF���v�81�b�Z&A^&Gcf��l M�������a=����?L,� �������>�]~P�it2�V��,;�A��$ޑ��%��{j~i�����I޲��}���z�����'z�I�3�+\�ڽb�un��h�F�������7 7�m��w[�����a��1]�����>H�x����ϳ
���v^;��gAh���p�Ϊ7��[MQ�h� �-o��_}�К)$��F6$��|����>e���4_z�\�E�h�*���ue�/_
�Z�eo�\Y��c�N'�v�'C� x�Nz�Jm�㦴��Z��jԝ活U��;ql�	��ŭj��	��M�?��(X �ny�����W�a�,��/5�i����`_<�w��"�����ߵE}'��:�Uiy��~;)y�ۋ�K�p�����ݣ����3��1b�xĲu��&��� ����e���]�5��F6�}Q��%�+@���f���x �qO��[�[9��U������[��3}��q����J\����$�$�E${s#��ָvx�\����;]�����3ÌWT͘�����{q��߇��[�]2���*�کb+Ufh|sB��=���Ñ���/��G�c
uQS��b����Kw��� �2���c�1�[�'��C�W�^\a�0�@ؑ�#�VoZ�v'�M:��$¯u9�}�Y瘞�̗I&�*��j�NkF����:�L�w\ז:"�k��۸(��g	��l/����{�Xѹs��)Q�5V�=t�z��6~�K,kz���������Y*������u����7��Y[$o�sI��@k>�0:�a�ޏ��ثZ*J�e��f:̐F\	`|��p���D6�Q�n��5kfq�,֜V��1�S�Ѽ�\v=��Ȭk] �jP6k�^�ٛ$��k]��x%�Ԑ@=�����h�$ol��5�;��A�(�~��e�ѣ��ݻYZ��I#6;;v�H���؂]6���#��%���U��������+9���%vKb8���Y#�L�ؒi�����<2�c^�
�ڳ4u�B��%���cG2I<�C��Έ�i��s��!��׎ͧSg��o;��w ^c�+J-�\f��2訵A�fM�]�4�Z�� ��2ɰ�8��� �[,W�Ke��b'�c#��c�q����|��SU8��,�^��DD@DDD@Va�|o�
�����Akߥ���ث��-�z����Q��]�����'������U7|}*�}���n��Pa&Ȉ.�����,��������)�S�6B�V�A��e�h�Z �a�@��^��u�"" """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1ˋ�M��1�vKOa�5��T4�f�+T�ガ�д9�Y�#kys.n�RX���9�%��}��sQ��1��l۞͈��6H��2�c{wi����n��:L�Ӗ�v����̬��z�"��7RƼ������.D� �������w�"�V[$�4	c���\��~D�7}���^K��&^���2vl0��$��wZ�3��l�6y<����d�:<�dqu�E��DC��ub8��qJû؝� 6�PJb��1���R˦h�`��q��p���� �O%w�j���M���9q�uwI��}q�]��DO�����Ʋ�h�EI_0/\�J��$ہ����߇���p�w �{Ii���~��=�_A��ϫ|d��{`ῑ� ���杼ʢ�+��j�U���4�N�9$�A�l[�2ۘ
3��[�!Nlxu8�U��u�/�=�m݀�n@�j�óm�I�r���w���wSj��>�,�67��)"kp��ݻ��r���OW�%���Ax�&�a�P��;\�۱;ە�An�dv:VӰT��)ܳV�,k�j�ap�6"F����=�u1�sn�d0�3�r�RK@ޤ�}�ݷwa�-S�h��^�۫�a��!jY�|�S��緫<d������ܗF���f��Yq�e�����.�em}Ak�E�,PCa����>@���g�k���� ]�`�"mF�~��1�d߈e�/�:�B�	1��N��ߋ}�岽KKEGP��j<�}�I������k�\a����}��s�U�v"Dܯv�xe�^e'��ˢ�6���ZO-�w$�4���	�E{�p�	�EYJ�xC�O�^�+[������q��&}�8Ϣ�{+[��������!�'� ��p�	�E;��3�^���!�'�'���~��.���>�׭�=��RzD�,{I w�1���ǐ�ߘ#�N{)W�����n�{S��k����w|{��v䂼qc����������a��$ޑ��ꕞ,d+1�8��s�>5����>�A��{j~i�����I޲��}���z�����'z�I�3�+[�R�o1P2�$���&xxk��v���Go����d��?ҵ�՛�f)�R�Α�� Ulm ���$n܆�s򠵧����v��,�+�"�� sI�` �$�)�-֯����Դ=;��o5��b�t���M�8�� %�?��@G}�[�_sE���DA�k���0q��c��$d��=���w��_��es����x٩�L}���&�&|}O	d��7--'pT�IZ�+������Z�ea��mFdll{^\��F�p��^�:H��-Q�q�2t;�\V���̳>V��0�g}��Z{F����dt��Ժ�tYJ8���T�q�����5�����۟j��S��fcL�Ο�b+�2c$�ٶ�h�Y����:V����[��ܳ�cո����%X�^JX�D)��^�� r���<Jg�]C��ZҴpϫ���p�5�̂(��iK�A���ۚ��;I���$r���!��O$�h��ׁ��1�RgS���ߩ3}˳ok����S\�z6�J�b-��ZZ�:)䋈N��{�-ը�������N���'5�m����>���F��6u.&�)KW�^�~�~��@��m� F�py���s#�p�j�J�f���׮����[$���n�Z��$�˞���ĺK.*\��ⴎm��q����pv<��ź��d,;H�ݐ�	�GTI%���\�\��w����(��ϛa�T�Y���&���y7n�wԽj�Xx�����U���խY���
��#�����r�;�_H�r^�����M{+��{����Ŝ��onD��L���Y#'`�I��˱kZ��ƶ���B�Ԫ�2�lă&���&��9�3���=��##�x�ˀ/xB�#��-L��Y=9��v6��vN�(�hm� �F�~s�w�+�r:WSV�$��c��q���2]G׊("�6ݤLI� ��w~�!������t.��Z��,�q���37����9� �w� �d����I/��7�~CnJl�� u�
MM�2��^Ȧ�]���f�;J�#�#/��,\w+�H���;�h�ih#r\O-�o�:���Lc&�6ȱb�ϒ�q����$o}#8ᓳ~@�䚏t&WPjK3��T��p�e�j���$�(e,�l���n�#�'n�zI�DW�����qeߵN*l����uK�Is��cs�@v�c��������W��o�k��ֆK.l-5���f��;(M�.��.�N�[�z��6e1R�](⛆�vE�v �8��;��v䗱ΖK�2'�'cg�>��\����4 �s��<�`UU�4p�yN'�lD�h:ǣ,�Y��j�b������$�07�ޝ��s��v�2xs�a8�CR�� ^�� ��`3�oiy۱N��� \�ݪ�E5'z;���/V)Y��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A���/c��c�3�� ������r�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ܴ��Oc>K�
^t���2��5>~��7�Y1%���47���O��{�ϒ���*���Fd��+�=���6�g�6g�� $p2F�����惿T���X�+'�f�#�75�#pA�#Ʈ��������.:�;��˘S��e��c��c;���80��F�n��Q�1���e�5cmX�j�4]����4F�܏ݭn6�P}��ū�:I�Z�+7����)� �Zǂk�����n69�^K��sV�:_�&����3�3fЖAB�S�������8�[�s��C[�]*7b���5��Ygs��њ�I�c��5� q��F�ݗ.��S�թ��Z%�W��r�O  �_@����O�ϵ|�L˪'d!��ڸ����݇c�\7�ޭ�� b���p�˻'��7����i �dxa!�q�~|�.]ӭ��cOk{�ҹ��q��-CM���'�r0��c�,���?�<|� ��!���,S����g��h���t�.-`'w84��'Ĭ�K��*y�=�^��i|6����|e���=a�5�wU?Jc�ä���I$�jT}��旗���䝚O�󃫦zU��m)^�7X˖lŅf|}Ǘ��	}�\6Y�����ڃ���r_���H��m|���7���kN�Y:��4as�յ�~Ŏ�w�s];�R��hc5�9j��Dr�f����%wU+�X��]��wn� �(����������=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$����f���f��c�b�z��.��n홻�]��l��g�Tc~�V���F����2o��n݇`�ߟ�����%����8mA��F(�C�������+m��h� �-Nh�t�S!i�)��b�q���q5�8���o���wߖ��_sE���E�A�j�:�Վ��E$��u�+�2H�p��p��a�f���f�:I�:�K�»! i���ּ9�cx����6�,p�ak�-��2i����E��B6[1K�i�sIo1�rA6�¨����3�f�q���.��Ӫ������w1�a#+����>bIf1t�5gK�k��u�et25���ih��!s��4-\��u@g�����e/�j��z���+�����`+��'��O洔�GSab�ԟr�
F(�s:ݛd�������@��[:�G{QK><��iY��z�mB`�xH=������sAԆ�ӵ�V{7���KD��Z^׽����&�#�ݡ�>"���4�K"�}<�2��7��`��#`w}� �v��o�c���2�k�a��ck�.�ۮ:�$f�p�2Y�h��nx^����Cb	��#�O��������>͂�����g%r�
���kR�6y K��b������IW)Z���5yD��V����b@s����Ngv��O-��q�3�x�� H+�>,%�C,���Hu��+��~nq%�= b��-�6z��3�G��}oU������z<|��S!V�mk0�uy36'�� �m��ӱ�U�����uguwd�;,�Ӣ�=\�� ��87����ŲiYoOJ[���2;!a�G��4Ms<�\OkC�� ����5Nw�舍DD@DD�������~�J�����R5��y� q����j��t������|��uc��������{��hݮ�7#��Wze���Jj�d��:���_�`q�d�i��b?\<j;9��tR�b��P�O��fN�|�[��1ɿa �g���^��t�8ߪw�?��'9lXN�09�U>.�r���e����ˡpd�c� ���� ��5�ia�Hi��ck�H�+H��$p�	�����ž��Zv���%��4lٽZ\V2[�Ҏ8șε'���f��6��ض���` �'��vY%���pp�:G�G"�����<�j�D���ОDEΑY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A���/c��c�3�� ������r�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ��v��N�ね3K^&���w��VH3����O�X��/a�\ �3v�	�j��Mj��m*ջ�dj2���=΁�T2c� wϑ���ͱ�ȃ�m�$�:�D� �_'=�DP^��!�!�����, |N��Fݫ��s����R�77S#�3�Y�<��ӎecX���Z�����v۞�ۣ�M�z���NxceG���wd�{9�������n�p�]�\�SV�BV�rx��}����s���5�h'� �,��îD� Ⱥa��V��l]Ź��>��qM�����������d����E��j�`�y,vI��Wau,�!#�/q��-%��"y����'��_�⣳�pj�D���,vS?[R�dRp�9��܎�kO���i�d􎦓��S�I�t��`p-�\؎�.>Ѷ�n{����t�R6�rm֝�K�8�2.tE����6 .��n;;J�����O�^�d����j�gO�W�'��Cr��u���*IF��u���)�S���'��$A�S���'���O�_�⤑n�O�_��e>���D�e>��m��u���*I`ҳ`�|Z�0���=�#�r�ǹ&�W{.0>���rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$����f����H�[wX���`-�w�yېې���[������G��ݘ�b�,h�`k�\Nٛ����M���LenX�]�vc3���	d�|}_X�Ƃ��=��V�W��|A�Z��6�͎����Y$�c[ָo��{�?ܶ����RȨ�Bɭp1Mv'樶JM/��X`04v���@�1=3Ѩ���G�R��^٣.�.�{�]|�y!ٰ���6֭��}�MJ���<��ы� ����ϑ#���ƴӒb��&c&=�_3�0��i;�^������U�U��	��8�q�^�n���N��g	ݜg}��I���ͧ����c���Z�l26F6b����< ���U����>_���G&.�s�jx�%2�!�KI��c s܇yB����^a�����nW�V�PC�c��n����z��Q�j�L��.�	�Y"�i��ց���n�w�%���|^��{���n�I����`�p� ���v��lWT�H;ϸ��{^�w��"�D�w��g�ʂ7hܫ4���Ɂff6Z��6G7�;�3b��p����jaj���ex8�'.'����\�O�f��e�5R """ ""6M�������T��������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���m8zϗO��$��e��pw`����oN���3�}@�OOd���]Z��������nf�e�)�+�`��xd4m޻�A���{\~����۶�����7��S�i�r�����c��,�W��C�q���جΏ�}��&f���{!�j�v��b(��tnw'��v�FSMÚ�Z����<P�4<E�pyo����L6�®E��p;�dn�f_)���ƿ��V��X�;��L'l���um��p�d��)�_e~����(��١R�a}'�ۦ��&dRC�]�F��=�������m�-���q�/�?��̎Z���M�b���mY$��:f� �6y&.�������}����u�/3m׹d�6G�]�\��3m�1���_k�Z� E��6���]�V��� t�kZæ(Ov��:��DT�uf>HD���\c!��s}�.�9��_���.�)�� -����������m�_����A��� -���_���.�+1a��_�����������D{_���.�)�� -���j��ç��s�x `���\�1�I�#���{�oH��[�}���z�����'zʧ�����
�~���(1'�����&���9���q@C�yX����������ߟ�i��3�+Pԗ+�Pѭ싫[yc�`Gc���8��k�4�"t��H%��uDm��%�9�y���|�w�GsC������!����j*��>A�7�|Oi<?��P�1k|֏��Y�{)U�+㵒��_�"�4�N�N�Ӿ	��W���waz(��݇Qq�.~���vU�Er��k>ŋ2�{�N7��1m����V��[:��=(gࣚ�H��J�rG��<�GY�۳��k��{����^�3�AJ'cv����x��;Is;�� �}��uڵ\N)�vڵr'��M�tSr|�l}��XfF�Cb�W�s^�$.m�m�g�}C5�쾰~��V���;�y�� �t��f�Tn[1>)�G����2�f;rގ'�ww d>` �E�+Q��e���3�pL�{������qI�y����J��r�ݪQU��b��O����F��;���=/_���`���2Թ��<�i"1P���Y�������G�5��M�]��[�v�uf�ZH�t+���k����@`���e��8c��8}�(�X��/����m쫫IzV8�J�5�H�k���� ��;-��	�N%�1�8T��""" """ """ """ """ ""�����W��|$��{^�(��_��]}yo���Ȩ��ҏ����U��ז�=\�%%�D^����[�UKSw��҃	^�{���g��AG��c�3�� ����������������������������������_�G�V���Ò��?tſU�_�}eh9�|9/�3�LA�i�{�ϒ���(}��^�s�|�R�l�0c�Ϩ�1��#q��fݝ�{�_�𰸞���^�v�0vZv?<�����G��Q�#EF�I dn��O٤n6�G����mf�MLōghFrX���m��tKx_��͠�� �ش@մsKd��Km�,E�K#|A�Qf�s���"�x�[-ܮ���2X�{�v��9ĶW�3���W�c����2�{lD���cC�H��A����\�����%�R]�H�ͳQ[�M�3�Cą�n�a����f���N�~�̴عe��[P5��V��k!ګ.�'�c7/&2<���uH,IA�&���K ��r��#2<m�Z�cncm��GT`*b$�2y�!e��tF3,n �|Cq��yPh���G�[,����5�b���eH�`���1I��]�', ���iY5�����ϨmZ�c��rܐ0�Ȗ�Y�F��%�f��ˠ>���QMW�FO֊\�D$���v$���LΛ�8���e�Y�#���ld6N!� ��(4L/��#]��D5%�8��W�7�c��>V�'DG}�����l��{��Ӳ_eX�t�wW����1�`ݜN��Z�s����Mg��;�f'��;�f �E����Y�����Y�$�F}�c�b}�c�b	4Q�k��Ř�k��Ř�Mg��;�f'��;�V|�$��{�oH��u*5�B���Bc�ߐ;��r�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J����nZ	�O��V�S 7m�+>(#��M�����7�O�ARu}������ݹr��T�$<E�S8�i��y�9��U��-tm-=��H갿��6����v+���2�jB\\baq�<<���R�66����b��fLʆDؚƆ���U�� DDD@DDD@DDD@DDD@DDD@DDD@Va�|o�
�����Akߥ���ث��-�z����Q��]�����'������U7|}*�}���n��Pa""��uX����H(�w��|FzܤY��H���s��r_�g�􏬭;�%��~�6\V��ߐ5��ϗ�P��0�F�VW��J+KR܌�f9=��b���]���~rſY���È�
�I�5�:8�mױo,,>S��5�;��u�~���� �hiX��=�u�嬺Č-ۄ:&F[�������Td`p���o"����}��&�F�Y7�F��Ӄ�k	y���y߾pi C�+����v�9[�Xn2:QF�@�z�oϿ<Lh����u�����������4���ز]��,��݀�/in��~�G%]*J�]q��kيW�������؎�=�=/�b�)�=/�b�(5��=|W(�܈k+6��@�h�!��Wm�{N�-�,Oa�~+�Oa�~+�A���z_���S�z_���Pf"����}���}�������_E=����_Eb,?a�~+�Oa�~+�A���z_���S�z_���PR��e߷=� ���NcܓzG��W�V�m����9�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J$DA{���)��U���[��" """ """ """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1��k�k�7!e�r��V�1�Vq���y��ty��� /c?eg�Q�Ӽ�F����˓Qc^�Η�/k�,���q�ί�E��� *� HG�W5���z2�7q]Wc.K���8����o` 9���ץL���Y:���1J
t$FH0>W]�$w�"-k���`7#nӸ)f���Ԁ���������7��w-��s�4�a�}��*�A3��^���#����ix��"�j�~�ͨl
�K�Y4�0���6#`���w�����zgPj��L6�7��be�r�I.>��ug`�1'�><|��}��~��1 �R&���cc[�֍�@r@�_��M�a��wF�Y��&E���N`�~�ش5��ȃ��>̇Գ���!�4�r[�d�K��tUs�ޯ�wxn�m�km黤��ך+�h��S��^��|��]�"������~��O5���SBT�r�:Ok��^�M��c�A$�pۘs�q27YYΉ�~� ��; D�����CD���pc7�����e�=�����qe`�Xmo$r��#����%��b�.`���@��OQkZ>�
)\9;�`���#E��J����p�ۂB�2�?��ͳ1&��;(�6Ѭ�0DF!�o���G%w�V��?Nc�%t� �G0�\����9 ֤��:0������9����2;z�tN���{�hoz��; H�����nW'z�F[Ӳ[�sAk��u��6�hf�4���m�.�/G�zl,#���&�Zڴ�`G ��ȑ��VLzC�c*���9��� ���p�4y A�*t�����:�2�
9�̓A3c�'�J�K7sxC��vqܭ�/�m�#���?�תD�S�G1�}Í�?��v���7a��-��G��7�k[WN��F��6k�o��<]�o/���]��c����ڥT�����o�!�-��4��/گ��y��h-a��Yy���%��y�pj	����^���a	��&�Z8]{�-K�K����ʠogk�vs߬t}�-�fi������1tCg��p9�vl[��9(�a�&X�7mW����m�#��jخ��|�\��t=����R���}zx�q�lG���6g�<r4��9��vp=�|\�r��i6�V��kT�V�d��[N�m��w�y��" .7��$ޑ��싍�=�7�}`���>����=AUO����eS���S�L�U?�N����g�U�r� J���<�I��4_z�d�ނ����/�=H.�"" """ """ """ """ """ """ """ +0�I�7�yY��M�� ���ҏ����U��ז�=\��^�(��_��]}yo���ȂR_tE�*����T���U7|}(0��w��|Fzܤ~;�V>#=nR��������������������������������,��_�}eh9�|9/�3�L[�_�G�V���Ò��?t����o�Ή4�O���e��]a�mkz�#�~�K��{�Pt��^^z8�bX�оśvk�A^6�����o�?�+�}�rI_��m��u�oV������D����_=���F"�8=�d���-gLm �&�u,>(�ql6��s����l�>�f[�4��r��7��N=c>�=e�n��߱��x�M�~�y��� ���t�cRt&��.�����;��H�1��˹ i!må�^>Yk���Ӷ�ԖW���	K�T_�K���۸P�ث�٫~��`��H��e�X�����#7n� F�m�5�j�u>B�+/�y<�y*#�mF�jкG��q.��l��.ݗ�^ջB��_�MS�H��l����Y�s��o#�M,�cs0��v�~������s���� �����N���-<fA�lF�ީ��K��\6<$�vߴ.{O�u�R�6ݑmɦy�#�U˛;�n[eѵ�?�O  � 8yn7[~���j�&v�tƄ  �����R{ym÷�y/Q�����/�ԃK��1�o����C�Y��sx; Y�>ɼ���o�2X���R�6�mb��؍�{ZC��ؒ������������l4{�<mgn��Y]7�hpm� �-礏��N�.�liL$p�Kn+��6�C����vn\��nOc�S���-��T��k1�q�ə�G���:�bsZK��F<�jVˏ�C�[��:v�1���<N6��W��s�s9v���s���1�j��5�P��*ۂ8��"�����wF�$��bӻ�ztGؑ���=	sٹ�3��a�5����X�#��o/�Zҝ%�qz�<f�N����'v��x��n�p����-Kӎ��#�6+Mq^��呸��c$;�k\	s�At+�<R�b��*�ߐ�Յ*�l K�xk���؟ �7$�����7g�k>��H�9⭇L�<����2F��;lT�g�Sѷb͙�w%���d�&������hؒ�6 nvS��y��_�S�}�f�:�Ym����$�=����i9�f��=����7`e��s���ᑥ��- ��p[���)[RW��Y��(h�4@N
���1��/m�����c����JL��1�F�^W���8�7k�� Gn�G��:�#-nA�mF$%�[����.p�/�O	;��u�n�#��3K>j��P<�G���!�I/���l@+m�]�N�qW[u����1���6Y9=��K6��v��x;�����cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���L;'J���En���f�X�9�G�v��y�Cw� _���^���� �\�2��O(�u[���Q��fq��RX���Yώh�`��s}�p�v�ٷ4��<Y��C/N� vu���L�[/V~�i#��o�Ƶ�j=��n���-\��E8��4�n���7�"��;��G��qZ���J�F㢹�;��U�����$=�!��p��9s��+�c�>��� ��3N�;Y,krqeE�;��y�CkE\Wcl�����lCO2p�Z�� H�[S���IA�κ�l�֍�A�bp�3�n�w=¢I�#��\�ےv�J䚃��댃�������Z�!]��'�Źy�JA�>٧�m��c���P�T�0٧A�����3�ͪ��:����̖:#���o�l� �t��c�߿I�v��/�pu�j�&<�\ �2k/n�r���/�Y�܆���FɊ����H��K��e+W�+k��Ŷ�^��1�s��xx����{<h:}�i������!nT�ر�1��n�ý��G=��[pݭ�%�V	#{{�7r�:��mN�k�oc)��L�vI�-��OT�����_�{��������t����&=�g�$-��#atm������������	=���rt�c�85��y Qc�&[�Ym������� �H$�a�n����L�JnP��9#�y[d���5�}�}߃�n��簅��=M���U�_"t�*Bg[t��X��"��9�!��GP}��Aq������Tbngf�hW�q͊I"��E�1���ηb�;m�\��Z{Wb�Yء��d:�{3ъ�=v9�f�0�9�"i�����v�!����4��0c�w3�3)�����q�0�� ��r'}��a�뽠""�y�rM�X.ȸ�cܓzG�:�3�mO�3�T��;�U8Ͻ�?4�PUS�?��YA�?��[W'����h)����T�_sE��FI���*N�����Ԃ�" """ """ """ """ """ """ """ ""�����W��|$��{^�(��_��]}yo���Ȩ��ҏ����U��ז�=\�%%�D^����[�UKSw��҃	^�{���g��AG��c�3�� ����������������������������������_�G�V���Ò��?tſU�_�}eh9�|9/�3�LA.�T1��L����C�\��2c�>��A#b'�� �7�G��n�*�(�-[p�f���E+C��+;m���lE�?"������7���Ɩ�e���<��sK�{�]ހ?� 9)^<K������H�0��>9�Q���#����XVz@��g6����2��`�-���Й�ٖH�1�q�
і�v����;oM���}�֡������?UnW���$�[���F����fa=��=5jgM�T1�c����� ��A�� �l�	���m�w]�l
�=*�+��7�����m�m�uۏ�ַ���[w��wk��w1��/�+>B�H���e��v2�d2k���6���n�n|G��{d��V�Gm�0I`�nN痤�s`�:�S��#U^�7���d*��C䉌Ŵc�9�3�{��a�P���<Ί�x�@&��Pf1»�H�摷qp�<�o%��!���@#}�})�N�\B�L���?b�;H1�{"��<Ld���k+�\䞳��<js�~���,�8)ER�q���J�O���ֳ�\��m��A��	��؝K��Z���4�P��25����9ƽh�tqE��,q<��gbw�e���Xg#�3ج}93Y��b�N�d2ֱ1of.s��4q���/j6A��G�8B��$t���Z�/V���Xz�9�e�2<�fXH8 ֶ>-�>?��tը-j|�+!�c&Ȇ؜I {*֣.���|]i�'��܈!�v^�,&Df0�/�ub�x��~&�m� U������=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J$DA{���)��U���[��" """ """ """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1t��ˈ���ͯf�5���A�Ж�c��د�C�v��C� ��� �Li�p��&&j�I#����(?Ϣ�\�a�&#n*r�%bY��\&�5���aϒΏM���N�3�f5�sPB�>^�R���g�N��}��֘5JR�W}>��:�m��<-ݽ�a�W$�be./�Q�΍�.cN>v�6�x�gqW�>�w��蠎L �RqJ���:��uLⅾ ÷z<�Zf���e���h�'}�r	���r��R��_�,�(i��}5�X������8h�w3#h�rx���y�W���ӽϒ�)���F�\$-2����o�q�?�}�*� �g�A�����q{���*���'}�`۽��{#���&�k��ܖDrX��s�؞�!�U� Ϣ��_�,�(0���g�+T���&4�����^~�j��Z4+���㉍=fż|����o۱>U%�U� Ϣ��_�,�(1lQ��|�*Һx��W=�&H��o���ܻ9��KN�1�,����ailP����Ð�0(h�)N��}�*� �g�A�Rւ&G�dlhkZ�  v }��Y􂧸���E;���Y�PU�P��H'uC�V} ��*� �g�N��}P��H.A�;ԛ�>�]w����Er�ڤޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���d�����ng1�A�BǾ�&B��6.�x�Ttc�>��q�_���!�Z$��s	> {	�-�����t�[��+MN8�F�5�, �j�Ki,N�����чB�!��9>R|���&�bbw�G<��,LLn��q�ֻ���N��4�l����u�Ů�>&�͉��yU��1C���*��ͨ�䅗������8�"��;��ndm�[/I�/�2�o'��T���O,����fI��ů��s�%b���M��kT|�81��|�;@�o>З;o�t�6��"������9��ej~���4����̜U�H��~��_�����<x���X��솩���kt�F�;=xn_��p�LՐ�Av��l��� c�wZGq�3����b�j[�7Ǿ�A����N�a�RY�-��k>�B�禡+_���~�pF������LF�"3�� �f�\��93���7�����T����OǹѺIe�9�;��'��%�za�{*T������ʗjL��D�I�o��*���=�EO?��3��)kQE{�0Y����0i�gM�NO/6C%��A>r�Svi��Ya��&D����ے|cȭ؈����� *�V���#��� 	~�,<����Ѷq��S2�Lꍐ�������m��?@��_��P��dkѲ�$��{Z�w	�$���؞~E��	�U�n��[�r_}�,c%���\Xى�8� �����KOk�3�sg0C4$R�+:�:�	�{�" �*�Ɵvwz��V�z7��]`/W����DD@DDD@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ���%��"����_�b��H�� ;U/��k�=�~\���X�.Gr�S��c����ii؍���G��W���o���o5�G5�E��J���,�et9��1���88yzW�k��꽋�錰6�BZ�Be���$kx��s��i�����=[2(���ꊓY��e�!����8da��؏�� �EFT�'Oݼ�]��l��⒬̍��\$c^����v�vMڧ�ħ�jE���V�c�ީ/]V�M�)6#����y�eq��U�LOEh�����T3
�Q�<g����iblc�`C-��Y�$���>NC�{��a�И�F�G�I��XDD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%�� T~�����,_P)��t�S&���hZ�B1Y
NeR8�,�A��H��7��[�֗KH�*�<U�c.�`V������0�uo=�����ݿ>]��]ԗ������o��eDV��ű����@�oX#��E7��b0��WVf��/V�>�t��U~���n��Ȣm�9��xw�o�����-��+2���d-��̲��0�q��7�b9��(����`l2�w�~ܭ��c)ݵ=:���!�$,h{�o|G?���f�)��H�1�WG4�ؼ�3P��4��dl�q��Q�{ k˽�h>?Ql~��GiN��ۭ���|�,��%�CMkvw6��.q�ɣm�]�`���}����}�ވ�^�w�g�j�/ӉѰMDG�9�<N`g1˼X�s����I��+!�/��W"`�y�n/�-��x<�«7��ϪcODDS����5)��[&&��2��"��-s��ͷ�4s�~~+��e��q�2�,}\�Xy#�P{��S,m#r�{�s|e�s�}���9����#��{.,c�F��� *��c ��e�x剆]מb\;I�;ٺ�24*�f'!.idߩ��&�w<�H���aR���C$W18;�15nӰ�qۭ��	���l}�7��p��Ej�S��`���CYm�@��~ffb�6""e�����G�oˉ�˧r\X{�|v�rıp��Oѐ|[쥛��k�E�X{r�!�2۟(\=�kNȚ;�\<lo܎�Ǻ��!{�q�ڟQ��U�;6^�gh����=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J$DA{���)��U���[��" """ """ """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1�=�b�K�
A݊?N{����/���A��Z�63W��$�ɩKCwJٚ��Y�T��ڢ�?%#f?	��{��3J��Gk���cd.÷b7N�o��m�۞�zn�ӌ9*��V�_4�[8iwA�|��Gڑv�{���R=�~�p��e��W��b3ڃ�2�*���<�l�Jh���w~㗍u�䀹��X\�M<#q�CR��:� ��h'�V��5�1�J4�Q11=#�/U!�/C�\�稼�U���CʜCʁ��q�	�q*� �e��p�@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%�� T~�����,_P)�C׺��+9��Z�$XC^�kq���c�o(���?Z��sX/c13Q�'�mX.��Wɽ�xZ������%�5���q���˵���'as\�󀱲�'��A��X��Ml|L��k]�ּ�w0���k����]��Vh�9��;7sD��5�4����IN�����Z׻�]��y�'J���F3�f@⌂Bl�}�g�nݹ���F�v�-�����#����ܙc~�o������W~а���.�@^�2qq;��,��87����x��n[�M�]0��Nw��3�[�2X�ѭ'��bZG>B��m�x�g�쵼ĺ�c����xq�fLD�q��s�|��#�HCK�ϔn�y�M7Э\^RŻ�Yb2#�+��d�h9������\�[^����n���	gtB	\ǹ�t`� im����3�V߷E_�������]+ޚl�1����YfK1��1�Y��~q�����9���3�,���ߏ���	j�la��k`|� ��˰��[��?#���\vY��c�����.d�w�wr�l�6�G�J�Vlu�]��d�����[�瓻�ӷ2Fܕw�GHN��˟��)��W�[ަ��RI�4lh�v��9� ���q���CZ�uy1vb�/^��e�3?���"�͙��M�3˴*�kte����<"h�c+����c;4�.��,��~&b�� |WdȰ�V�5���m��&�_�Jb�����KW�������c�~�;�?%bf�@����� H9)j]'g2yc������nĳ���=NΉ�hw>�n`lZ{Gn���n?-K���\�αr"	H�q������*1��1R�`��1�X4��G���q�9ė�G���ߵ�D[�����Dt����;��N,p������&ys�Oa�T�����bg�GU�P�5���3��9d��2=���ŷ�m���NG�m(蘡h�0�+��uL�Z�x�Cۃ�n��Y�9SPԣF���iC]�dh���� ���~7��b�S<�E�c��i:�"�����zB����&0v4 ���DD���=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�����)~�t=��~O_�"��ķP@A �����iG��Ēh�$��A�KSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%�����Ӟ��%����w%�'��0�f23^�+�dy�:'@=�=s��x��1�)�mimd��:�b�=Pp.|3=�o2���'̶�I�����UoɎ�Qd�G3׃�m �Ll;��P�>�q�,.�3���"~��qXi$�� ���@�i�x�������3;��D��t�&S�b�B:��^`�dM����^������ݖ��V��k]S)R:7d�f:�{�l�hr{� �Ϻ�ԝc5M�ܞ]��W�X� ��8g�Ƿp��[.�ӱi�|�b��6K3Y.x �$�y�]�\����������Lv���^�gc�	�^�DD@DD��ר���"" .7��$ޑ��싍�=�7�}`���>����=AUO����eS���S�L�U?�N����g�U�r� J���<�I��4_z�d�ނ����/�=H.�"" """ """ """ """ """ """ """ +0�I�7�yY��M�� �s��oSV��q���o��خi�ϧ���/��f��7b�kߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%�� B�Ӟ��%�� Pj�X�����UjM.B+��-�W�p�nOY� E��󋧒���j(2�ϹF���7kz�N�`H'�n���.{	���t���b'A������^�ly�� �@�:&��%\��a�ڥm��LAatqw�5��'��w2馛UDoN9~�*��MS���6x�L�_�CB�vs���#�AK	o~	$��O�*�����:��&���L��;�p���@<$�O=�����g���s5YEjй��)	;1�m���ǒ�gA�*�
��A�qSo��g��6Bx��m�s�U���W%f�G�-��JG�ԙ):hq����0�(��7vxM�#ī���#� f<?"��q-����枳}�G�#o�u��z:����d`�f��F����k�nmcG1�e���.�[�E�*w8�����o����~+Uc���OF����oFy�N�c�{;�a�qH�A���sc����8�	]V��tɶ�M�ȸ�����ɍ�����Fxe͑��F��4���<��V��^8�ܱ���^�c���8ٞ"�".g`����������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�ܰ4��_�b��H�G�)i��מ;6�Zl���HL�3n7m�M�Aa��'z�Z�S�kc!e�����7F$k�2�zZG�Et�������E��J�Z��[��p�Z\洰����Gůe4F��O�Yb8��CW?4nkCY���o�x�;ǟ馊&�̸��r*�������u<ZxL��$���'0�������r�ۚ����݃	,rI��{�T��nZǽ��;�ܴ�5Dڅڔ�^9dH�<�P	�ñ��xv�ڰΓ�V�ؼ!�I��]�㥏��_�F#�ۂz�Om�V�v���� p�]�iu�9(k;s#^����'�|�0��y�]�;l՗~	Z�c���;z;�U�c⯋lx�q��ƹ���l���o��Xn��v[�D�)�΋���@c�$�,o���8I�Ao��UQM4�%����V&1�.��{�oH��vE����>�A��{j~i�����I޲��}���z�����'z�I�3�*ڹ?��[AL�ނ����/�=J2O�ARu}���Q�|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*����H���;�V>#=nR
?���)D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDj�/�>�������-����#�+A����~q��b�N{����/���Ӟ��%�� Pxv�v���V���M5)L0Yx�e�����N�#9m����^1�ڶ+W�G�[��ւL���Fɞ]��;����]�ވ��w暦0�`��a���l�F�{&lw���U�����+C{H��ٰ*��e���=��܊�?*�W}vB`6�n������G�;�GXv�7*�Asތ��s��+�Y��w�ꡘ0ꐿf�����~����Ж5S�VW�N��DP�DDD@DDD@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%�� T~�����,_P)��>�E���Ee��l� �
�Ձυ�C��ݜ���䴞���.W��ږ<; �Z�<DǿY�{8���3ǲ��]�b}����Nm�MGq�I���Xs��������Z<Am�i�K�n�M3��}W�m�V��Z6lŀ�j}W04ֈ�g7��m����� �r�1�}�cDͩ-_��1��6et�F��>-�=��̲z;ԙ�֭��6�L�~�mA̍^�nds�����@�nfl�3����U1]B:�C3�&2W�����7>=��y�Io/u�)�;�x����,������s{��"�=%g��ZlEG�f��o)_�c�cjF��8�����o�"v;�E���w�i�0�� v�u�`�;��IlV�V�y����ax�qunq{��;q���ﺁҝ*g(�
��v�#V�I�^�ٷ�o�Vw�@i��."v�ڣ�\�N�DK�l���8�2��
.��tX+�ݍ��D-����.�a;l6Ue��X��]�_d;�#&��V�P���w�7p��~[�3�ޜ&u�4�]��̽�p���CG��J�E���-��o�@��6l����'��E�����I5VC^�:ח��m���E�^�8��Uji��j/�s�7DDX�DD@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%�� ����_�b��H�5�CS!V+���'U3C���ӷ��V.gI���I���nH�k#w y<��أ5&��M�|Wt�0���d�x��3 {N�B���B����ނ����fV6�-t���C��ʵ�k�a�U�7�f9�wi�c���P�>h�w{�# w� 6�/)�]��Fe����nŌqܴy��=ҴW���Jӥx���k-�h���8�����W�:C���$�JCJLov�쁍.wZ�m�v���
xw"'(���b!�C��G>q�5��������^Y���sCwPO�W{Ga24�T���-zM�g(��#�6 m�Z��m�	�P���ͷ4Nf�,�1�M�DN��C�aGҜԳ��~F�v���0�|�,��cOx	����a
�;��������i|Ll,n>��m��sv�O�6��h:�D=A�,lu��mZwh`y�"�4��kl�Z���Tb��Y+�n\���@��޿�a��R�����W�b(����G0,2̐I�ge3n�1��D\�\�c��c�j[9;�d�J&b���q=�qw��m��s�my}+��Cy
�m}��6�`�b� �����O�����<v��gH�F:6M����|�+g�g]u�3=QE�GTX�xƜv� ƒi���ZXx<��#�ռF�ܖN���H	v��hٌ�9�|e����ۯ  ��-7c�R"(\DDD@\o1�I�#���{�oH��[�}���z�����'zʧ�����
�~���(1'����j����m2x7z
���h� �(�<�I��4_z�]DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@Va�|o�
�����Akߥ���ث��-�z����Q��]�����'������U7|}*�}���n��Pa""��uX����H(�w��|FzܤY��H���s��r_�g�􏬭;�%��~�7=9�{�X��R�Q�s��/�}@�܃]�Z"����NE�2���.��.�����isO��b�>����1dnb����8��<���&���vŻ��k�_��"��p�e+رR�o�e�F��V�������~SY�f�bnQm;��AnQ�k����U����9-��M11��<*��f9��Ѷ2#b�x�u���Hن��h��v`���U�:?��r-շd��L�奲���w�����v��d^�U�z�LE֊��=��=����fn(Ϝ?̱0]$brձb����;(������48�qh'cϵ3st�����4(����X%�����;i"|�f�p���w�f��;4���0�_V����h%�nn��m̕��k^��c�R�u�b����H�v���F��F�>[Z�6^L[r��o����7�$	�f�",宻�����~s%���]y}~��6��i�0��6#b �+��Q���3Y	�HP��d�<�wX�\\�Iߞ�a�k<.��Xqy�K�l{�I��Gc��;)�J&�q�eh�ny�5��f�O��m��r�{�]��ll�6��O����6^��s9���� DE��������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�
�Ӟ��%�� N�5�e���th������q���lS�GI (��L�]oo-����w(ש#g�����$�$l�o��x�0���j�&d/��ck�v^+��1����@�]�SahЧfHVO]-�_+� ��=��p<��D�ˬ��k��ڷ^��L��cck���A>ԓ��`�&K3S*�R�B��-$��پݥ[�����~�y����44��9���<$G��~դ]�Lr�ʫ6��}\��DW�bp�j�Kqr�Γ���!˳�.��ɵѦJ͙+�=vb�j��M���N��F�����F�t{7#��\<Moz��;Cҭc335;���l=d�qlG|ǖ8s�9�$]��6m��D����-ݤj֭���c�i!���N� {����{����uտV�Z�-ӻ�����DDD@DDD@\o1�I�#���{�oH��[�}���z�����'zʧ�����
�~���(1'����j����m2x7z
���h� �(�<�I��4_z�]DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@Va�|o�
�����Akߥ���ث��-�z����Q��]�����'������U7|}*�}���n��Pa""��uX����H(�w��|FzܤY��H���s��r_�g�􏬭;�%��~�7=9�{�X��Y��Xs��/�}@�
U�.���l� F�V1�`K8����1�Rl� $ÛI�{��z�Aō����C]߰�-��H#~D�ۚܯeh�8;��x��������C$d�k��摸 �[qj���G7
����jz�M\�hK8�������z�,��lF�8�� m��.���:5��b��J�{�ś�*U��G<�u[����� ������%sK���m��A��¹�SE��Ev)��Ƣ��!��;2/��dV�p2��[��c��%�v����8���E��0Z��(i�q��<NO��k�!�r��{�r�;lƢ��S�����
3U�#L��/���f3䣙�d��+�������� k���QL������b��mZ���mÝ���T�\8B�˛��ѥ�|<��y����(�����0�nN��`O�+�Cp�t�E��z���������=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J$DA{���)��U���[��" """ """ """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1�=�b�K�
@�T~�����,_P)������@�1��R�Hjd7�~~�=���o��cɷ�D5ڗG\ӺB+n�E�h#e1���	p��Yc��۱vW1���!��W盗x{�]�O%�i;�f�vn��E7b)�f9C��335D�Θ920ˌ��z�y,~PI$�lo����sո�9��u���#7w!R_drS]�p��>��c�`8�hs�ſy�ڻX�$��	�s�9�ڝ�xV� 8C���W��U9�T�O4�"�4��Q�nd��r/�3'�nI��\�l7�D?ǿg�ei鵃�U��~J�Z��6 �c��v���>���>�ؘ͸X�l;�{��c7#�#�h�8�����5��n�/u]]<�-�b;��dQ7���O�F�����}:2��cu1+e���Yg��z{\�q�&6�����Tw$%�wT�'{c�7>��7�""i�:��3����::�!���e#5��k_+�&Ӷqh���eG��cl��^�PR}��U�=�J[3va��{8�j�De�\�}�۟f�%����5Br�s������pB��L�&6+�1SZ�;6��\��̇#b��Z:��@i�@�;V�n�����8S��6.7H�#˜����{I%IŅsT�=6�i�"��QQ�������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�
�Ӟ��%�� Ps���-J{y����vI#��;����'��@�wo.k�H9�lN#S��^�K�]���퓬�Mv�u�,b*Z�T�Iʬ�8d�������*�kC;e�H�}i"�U߲I6y~� � �ws;�馺1�tq�n�骙�.A��X�8l��ֻ+p��v+9Ί�k�����Ͼ�K��uY�����.t���ek8]ö�!�4{��l�������Cf����Ga�|�}�s��˳n[/!��OW��v<s<!�=�MgV��pgz��x��j��tڽLb*Dh}}��w�����[r�$s�[�֖�p9��<��k6��8"v�nZ�7Q71�i�wW7rί�����v���t�v��bf�-Z��Ju;�	<���� k~e�t�=���o[�����n��~=�qm��+�&q&�Ɉ��s�IY����� ��X���VW��Ogr@�zƞ]��5�iސ�f5k���Y��&���F�0@}2���)�h<#��X�i�:�Uk����k������ʝ;����gr�I��r0�1�"a�w 9۟'�SUv�&"M������M�M׫��������������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�y(�9�{�X��RA��A���q8,GsGr��|���8�1�8Z�I.��>�VC�
�L`��W�K+���$qɻ#ٲ;�����l<{�)�I�]��c�5nɎ�Rl��b65��']ȂX��![�CRu|,�=��6j)�v�B���\������[���e�1w3�� :K�]���خ���F���\��8�;�B׳=#e��Y벥L9�IJ<��$���6w�xi� s��n��G!�����Y�ڬ�Fq���1ż��;�죛�d������lѓ��k������Ȓ{��A>u16�bp�Qzbc,lgIP
Q3$Ɯ���H�)��������I�y�Q9~��ŧ�d�X|�@W�(ٻ�L��#�k��G�'gs��wE,���6�Y/��Z�$u�$�S��&���at��� �d?���ǔ�mI-�c�L#c\ޮ^��v����[�J�,�53~c�zoӵ2�h�l6h(s�ZZe�3$����Z�x�wiį[�.0L�K���������b��1J�vk��a��	ݡS���6L�fBFV��C勹�$I3�[�.s�ߴ�9,܏F52Qe�s�d)Ө� �[]�{H�3��W��Jc�J�#S�\��iס&�	*�8X2GF�x��߉������om;�6�GƮA��ȱM�o�s8Z޴���08�8�w�o��&����n��D~�DY�q�ǹ&�d\o1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ҭ���g�U�����*N�����ԣ$�n�'W��|A�AuY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A���/c��c�3�� ������r�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ����_�b��H��:v��ϒ��Բ](�����:~�8�9��+$�i}�	�v�F�f����O{��A�"�u������/kf��Ø�?�k���lQ���y�$@k�'�z�:��Zy#5co��?r�Z%cek��@ {xdg=��pF��W��͗����������������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nZ{��3�}@�{ZkT^�1�k��U�-p �^��ԍ�i:���һw�����q;Μ����,_P)=��>�)��?g+C��8����y���j�t�p��V8�a>��~�:/D:�G؜�I�Z���_r�+�����L1� ��������DD@DDD@DDD@DDD@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%��"����_�b��H�""" """ """ """ ""�y�rM�X.ȸ�cܓzG�:�3�mO�3�T��;�U8Ͻ�?4�PUS�?��YA�?��[W'����h)����T�_sE��FI���*N�����Ԃ�" """ """ """ """ """ """ """ ""�����W��|$��{^�(��_��]}yo���Ȩ��ҏ����U��ז�=\�%%�D^����[�UKSw��҃	^�{���g��AG��c�3�� ����������������������������������_�G�V���Ò��?tſU�_�}eh9�|9/�3�LA���{ؿ����Q�s��/�}@�Pq�ǹ&�d\o1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ҭ���g�U�����*N�����ԣ$�n�'W��|A�AuY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A���/c��c�3�� ������r�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ����_�b��H��9�{�X��R(��������������������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�Tv�����,_P)D@DDD@DDD@DDD@DDD@\o1�I�#���{�oH��[�}���z�����'zʧ�����
�~���(1'����j����m2x7z
���h� �(�<�I��4_z�]DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@Va�|o�
�����Akߥ���ث��-�z����Q��]�����'������U7|}*�}���n��Pa""��uX����H(�w��|FzܤY��H���s��r_�g�􏬭;�%��~�7=9�{�X��R*;N{����/��" """ """ """ """ .7��$ޑ��싍�=�7�}`���>����=AUO����eS���S�L�U?�N����g�U�r� J���<�I��4_z�d�ނ����/�=H.�"" """ """ """ """ """ """ """ +0�I�7�yY��M�� ���ҏ����U��ז�=\��^�(��_��]}yo���ȂR_tE�*����T���U7|}(0��w��|Fzܤ~;�V>#=nR��������������������������������,��_�}eh9�|9/�3�L[�_�G�V���Ò��?t�������,_P)�=�b�K�
E�{�oH��vE����>�A��{j~i�����I޲��}���z�����'z�I�3�*ڹ?��[AL�ނ����/�=J2O�ARu}���Q�|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*����H���;�V>#=nR
?���)D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDj�/�>�������-����#�+A����~q��b�N{����/���Ӟ��%��"���������������������=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J$DA{���)��U���[��" """ """ """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1�=�b�K�
EGi�{ؿ����@DDD@DDD@DDD@DDD@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%��"����_�b��H�""" """ """ """ ""�y�rM�X.ȸ�cܓzG�:�3�mO�3�T��;�U8Ͻ�?4�PUS�?��YA�?��[W'����h)����T�_sE��FI���*N�����Ԃ�" """ """ """ """ """ """ """ ""�����W��|$��{^�(��_��]}yo���Ȩ��ҏ����U��ז�=\�%%�D^����[�UKSw��҃	^�{���g��AG��c�3�� ����������������������������������_�G�V���Ò��?tſU�_�}eh9�|9/�3�LA���{ؿ����Q�s��/�}@�Pq�ǹ&�d\o1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ҭ���g�U�����*N�����ԣ$�n�'W��|A�AuY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A���/c��c�3�� ������r�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ����_�b��H��9�{�X��R(��������������������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�Tv�����,_P)D@DDD@DDD@DDD@DDD@\o1�I�#���{�oH��[�}���z�����'zʧ�����
�~���(1'����j����m2x7z
���h� �(�<�I��4_z�]DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@Va�|o�
�����Akߥ���ث��-�z����Q��]�����'������U7|}*�}���n��Pa""��uX����H(�w��|FzܤY��H���s��r_�g�􏬭;�%��~�7=9�{�X��R*;N{����/��" """ """ """ """ .7��$ޑ��싍�=�7�}`���>����=AUO����eS���S�L�U?�N����g�U�r� J���<�I��4_z�d�ނ����/�=H.�"" """ """ """ """ """ """ """ +0�I�7�yY��M�� ���ҏ����U��ז�=\��^�(��_��]}yo���ȂR_tE�*����T���U7|}(0��w��|Fzܤ~;�V>#=nR��������������������������������,��_�}eh9�|9/�3�L[�_�G�V���Ò��?t�������,_P)�=�b�K�
E�{�oH��vE����>�A��{j~i�����I޲��}���z�����'z�I�3�*ڹ?��[AL�ނ����/�=J2O�ARu}���Q�|$������&���C���G�r�v*�{��|���EE�~�~G/�b���������A)/�"�M��J�_tE�*����H���;�V>#=nR
?���)D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDj�/�>�������-����#�+A����~q��b�N{����/���Ӟ��%��"���������������������=�7�}`�"�y�rM�X �xϽ�?4�PUS�?��YT�>����=AUO����e$���m\��?ҭ��O�ARu}���'�w��:���R���������������������������������
�>o��^Va�|o�!�{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�U/�"�M��J$DA{���)��U���[��" """ """ """ """ """ """ """ ""5|�YZw�K����W�~�����}��8��1�=�b�K�
EGi�{ؿ����@DDD@DDD@DDD@DDD@DD����>�]�q�ǹ&�u�g�ڟ�g�*���w��q�{j~i�����I޲�� J��O��V�S'�w��:���R�����T�_sE���D@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDf	7��  �+0�I�7����Q��]�����'��Qkߥ���ث��-�z��JKSw��Ҫ��z
��o�" ���U���[����{���g��A��􏬭;�%��~�~��H���s��r_�gsӞ��%��"����_�b��H�""" """ """ """ ""�y�rM�X.ȸ�cܓzG�:�3�mO�3�T��;�U8Ͻ�?4�PUS�?��YA�?��[W'����h)����T�_sE��FI���*N�����Ԃ�" """ """ """ """ """ """ """ ""�����W��|$��{^�(��_��]}yo���Ȩ��ҏ����U��ז�=\�%%�D^����[�UKSw��҃	^�{���g��AG��c�3�� ����������������������������������_�G�V���Ò��?tſU�_�}eh9�|9/�3�LA���{ؿ����Q�s��/�}@�Pq�ǹ&�d\o1�I�#�o�����
�~���*�g�ڟ�g�*���w��ğ�?ҭ���g�U�����*N�����ԣ$�n�'W��|A�AuY��M��+��>o��=�~�~G/�b���������TZ��G�r�v*�{��|���D���/AT��-����D^����[�A���/c��c�3�� ������r�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDDAf���#�+A����~q��bߪ�/�>������� ����_�b��H��9�{�X��R(��������������������cܓzG��.7��$ޑ������S�L�U?�N��N3�mO�3�T��;�PbO��V���3�*�
d�n�'W��|A�Q�x7z
���h� � ������������������������������������&����f	7��  �׿J?#��WC�^[���r*-{���9~�t=��O_�"	I}���n��UR��/AT��-���DD�����r�Q��uX����H """ """ """ """ """ """ """ """ �W�~�����}��8��1o�|�YZw�K���nzs��/�}@�Tv�����,_P)D@DDD@DDD@DDD@DDD@\o1�I�#���{�oH��[�}���z�����'}b��}���z����c`6�� T�g�U���{ˉ#u�q3�P`I���*N�����ԭ���7<½:�5���d�"" """ """ """ """ """ """ """ +0�I�7�t����2w( �{���9~�t=��O_�"�׿J?#��WC�^[���r ���z
��o�_s������ZI۷��Y���)N�g�����U���[��ǆ�`��i$� w�o�U��"" """ """ """ """ """ """ """ �W�y����}��8��1t00l;>����~q��b�N{����/���Ӟ��%��"��������������������߮�m0F�YƂv� `\��R"�@s�����C�A�V��+׊/c*��`n��y�6�*���U_�O�o��$�֘�O���q�]��a{���{|��X������Wdh�Fb���rΪ�3��>]_�A�*��'�S�A�*��'�W(��:;�!�~�T��:;�!�~�U=�S�s������˫�!�?%U��� *��@?�Ui?ʹO�����;�2�����=C��T�ܵ?g?{��������<]_�O���U_�O�P߲�F��C��v�����oCջ��R0H�F�8����V7,]���L�[Qz���%)송��W����송��W�����)��?��O�L������ �`՛송��W����송��W�����)��?��O�L������ �o���U_�O���U_�O�/�L������ �>�2������ ��j�Ui?ʞ�j�Ui?ʰ���~/�?��F�ȉ��q���7:� d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���Od5䪿���Xl��W�;���#�j�2�d5䪿���T�'���s�Z֍�6N�}��ɑ�5~���Q6~��>7��c�Z@k�#�H<���֡���R�QW|C���I%��<�_|����s{��L;���[��?	C���A���e�G'k�#���g�=޷ ��CP�J��I�T�CP�J��I�U��ɑ�5~���>�2?��w� ��CP�J��I�T�CP�J��I�U��ɑ�5~���>�2?��w� ���A�*��'�W��j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʞ�j�Ui?ʰ��2?��w�'�&G����d��j�Ui?ʵ��+��=��G��7��ַ�o2�:�#�j�2���]���߇���۹A���{ؿ����Q�s��/�}@�Pq���f�d\o/�I�#�1�|�X� ����X�)n�5� ��տ��o�TwF��kk����bn7X�8w�p�}�M��V*���V3�_��#UU9�3����sK��7��Yټ�9q�r5�i�v���㑁�w"{ZA���:o��~���ێ��Y�p؊f�Hۮt��������vh�k���<�HZk?w#���ো��-��.��$i���A�y�㷯��&i�s�=��E4�Y���}��cm�R,��.OV�B�(���k����͸D�� ��9���zt�-i����d��K2�kC$y�^���6�5��lܹ�g�Y���Q5�YØl�M����� �6��_�ĿN:� �}�� �~���K� �G���� �W�7��|���9�iq٠��>e��/�u���k�/H�^ԵF�c�o�r�a�γv��:���O������Gg:HӚs,�nG&���\:�ȃ��2��-�y��^f�j9�Jq; �J�ᑎ�{y�y!�+���3�0X̠�Z��8Yg��N��-$��v���[�h��#P��V�q��Թ'Xp�᮪��,�o�ax��]�ݺ�|ǌ�ڢ�75]�ܭ(n�ju�ur�E�q�P��F]��m����d��3:QcZ/աZ�'c$�Y��ڭ�c2u��i"N0�C�G`�(|�� \���=lS
5�ʿ���������������������������������������������������������������������
� � �� �f�+� �?�� ������,_P)�=�b�K�
E���oH��vE����=a:s"��Ж���������5'�,�LȻ״��֩��:E۞����� 5��e�TH6�����eV��g�ch��=��_�5�C]LѦ�����~��ؕ�s_r��L����� ������ 4� @"� �?�澚��ڏ�m�� �J�D?ݴ6�?⽮��~_%�~����_6�z�Cz+�t�f�����K��ȃ��U�z�O;zK�-7��rM�����a�ܒ�������e�� �J�F?ݴ?��*8bg{�NL���Q���e�'� �q���~�~�tU����8Z�+IZx�W��sk�6 �����o��?��)�+u���� 2�u�/km
b���c�zz�vsAT�Eڧ>�����d�_��/���[�� &�� ����+u'���� �x_i�#���Og�ү�/�:��|��<������ҷQ�N�� �^��R�m�� �</�����Gg����Y}1�I��'T� ��|��+u���� ��������� �q���	�����K�~Y}1�<h~e��b{U�/sZǂ@�$�oR���V�=���� ����+u� v�� �������>aY=��I�����Z��d�2���.�+�� wQ� �������h� ��S��K�0}dl���.��e��?�Oc-~� 2�?ҷQ�M�� �O�[����C�� �O�/d|�~���U�e߽������e��?�\}����m��?�����?��=��}$���G�#�#�� i?�]� ��_�̞�Z��e���f�?���� ����a�Ρ� �)���G�Y=��I����Z��d�2���.�,5��8�$� }������L��>��:N����=�"��K8ݏ�[�`c;�~Y}�e��?�Oc-~� 2�_ҷQ�N��?��?�n��m�� ��m?d|¿Y=��I�����Z��d�2���.>��G����� �����h��S��O�0}d��'�˾�k�����_�̸���g��C�� �V[�[�d|����v�;v�{�J<1���1�G�>��8��_�e���� � �=�������~�L��	"������. � xr��+u!� v�� ���v_iOJ#�?I��ܫ�˿{k�����_�̸����h� ��W���{}�~��S�}�쏘G�Og��,�ﱖ� � �=����ˀ���Q��m�� ���Q��m�� ���/d|�~�6�O�~�2���'��� � �p�[�� &�� ����+u���� ���G�Y�*�����Z��d�2���.�+u���G�� ���:�?���x~������d�ӏ䏘D}$�~z\��˿�k�����_�̸�������W���P���@9݀���S�}�쏘#�'��� r,�� ��� � �=����ˁJ�F��>g� �����u�� �x_i�#�������Yw�c-~� 2{k��������m�� ���Q�N�� �Om?d|����� ���.��e��?�Oc-~� 2�?ҷQ��u�� �J�F?��?��)�m�쏘>�{?���e߽������e��?�\�V�?��>g� K��B͸�c۹�o�7>Ol���J?�>a1���&q*�����Z��d�2���.�+u�{���W�ҷQ��u�� ���?d|�>�{?���e�}������e��?�_?��Yj�/��h$4�;ڪ�����m�� �x_i�܏�O�F��w������Z��d�2���.~��G�:��� �?�f�?���� ���G�#�'�� i?�]���_�̞�Z��e�O�[������� �?�n���h��S��K�0}d�~z\��.��e��?�Oc-~� 2�'������S�V�=���� �������>`����u�?�]���_�̞�Z��e��n����� �T���2sn?�	��0v#�'���M����dlg�W���Z��d�2���. � ��P��=��{Z�0 �J��/sB��ر�͓��$����ciG)�>aj~��\鮩� ��о�Z��d�2���.>��G��m�� ���V�1��� �+x_i�#����� �O�}�2���'��� � �p/�[�����ߧ�S�V�>�c���S��O�0}d��'�˾�k�����_�̸���}���?O���V�=��6��� �<-�����Og��,�ﱖ� � �=����ˁJ�G�6��̟һQ��m�� �</�����Og��,�ﱖ� � �=����ˀ���Q������ �{�+u� wP���S��O�0}d��'�˾�k�����[�]� 2�C��c��@�?⾦�1�Z\6/hq��~���������=Q�;M��A5Ɔ���g1��_��_�̞�Z��e���Tӽ�����7+ZJ�!+	�mǡt5��_W��M��{ؿ����Q�s��/�}@�Pq�Ǹ��X]�q�ǹ'�XA֯{�o�W�~���]�d�5�'�5��a ����4�[����|�{�E�����g��S%g>�v��wi����"�.�k��(���q��/�{q�u�V暽������c��l�CoY[mg�v�k�tRfB�M#�������j�19e�nj�a5~�N)l���[nI%�G�Ҿ���F69���������5�s�O������$N��E�y�+x�����[6g{�ϟ��9�1���z�"�i'�?�3˟_�����.4�*�s�[��V��I�s��@-�5��ȭ�rN�#�mgE�g6_�g1�-�����C��I�����%}q_�k\�8� �8��>B���(>�yg����_$�W�kZ�_�-mmݙo3Şx����vG�:�����8�Q=g>X|S��Is=[F�He�Bܜ�D�9����}�=�$r ��iɲ50EO��6��]�N�;�r����X��z���5uL�)7�Z$n��vpy�7�#Y�����-m��jbb���Io��h�4�D�#9��c�>��z>H�ث6��`�q�-��BHlM p�w�� l<g��ːe�,2X��>�π���N�G�	�n����#X� ����� Rƥ�+��eu]WZ�b���b�;�F��ӳ�y��n��'oy礳��[�wzt�ˎuD� �>����H�T�Sז̳��	lO{"q������rU�;3����^�������	o<��}�~�k����^�"�I�q�2j�ܗv�ͻ\�7IN��[If�q���z��/N\��|���q���I3��;�5�p���O����'�i_�Z����r9+����9�-�߇�s��w����}��r�%:�v��	 0�?n-�ѷo1�W��3Tni�wk*C,�]a�LC�tM 9�{���	�na/m��vs7I4}������/�5>X� �|冖gcp�f:���W�>�w��j�KZgq�5�O�Ū&:��+�2oe�ؗF�3���I;y������(��)�u����Q��� �^���j�i��XX�nߵU���:���9ϧ?��7��m�U�J�C�!{:�=A���\��Fþ���t�!������\�6���e���ǵ=�y���?�Wjpܥ��۩3C��#Oak�� �B�����(�� ���O��6-E�n���>�Z��U�s�� �>����G�bיK�h��N27�9g{ח�	��ÿ�m��w��NX��e�TwouF���m�qwi�����G�������+V�÷]��X�A42����zGʝ���� �_)�uW�~��9]�1�<�����W�ZCwi,)$�i@I'r~�Ճ6BF�6Ul�u/��GPK#���;?��7=�r_SC� �^(�?q�����h�%b?�i��ǳVVu�bd���##y{X��=�\cx��;�WD��gMSq�yKϧ�;v/ݹ:\�y�8���I3��LM�#��HGU����^$"YZxO. ��Ge�����%�,��i��`g���Y�tm������g�"g���}��6��=�K� �s���������� ���m�ɦ�1?�>�~o��Ⱦ���Y�J�� p�7`��>�ȑ��}�vrQ'%=�S��fX}��+�qM��l�۞�x�ק�F�� 3�_�I����P��_�KJ��ϟ��s='�m�;nQ�&yDO�F'g�cϣ�����Q�[�[�%��������yao&�K�O��������Q����`m���!�܏j�ٿ������z��/t�$F2翱�<cr��e!_�?}��~k���4U٭h���V���Z�3U��=%mb�ƫOE6���ffyӏ�� ��1�+w���$�CIc߳wkH y7Z����a�v�E�]S��C4Mxs�yo���:���3UԔE�N����Ih��bX����!g���u� �� �[��̹N)�1�%ǥ�_h��8��b�.s1�~��ԙ����5/F��m��w��K.ݻp�c�M�qڶz�+�Ze�ǵ��\��.s]'=�$?辭?b5�����O�/�=�� �Q���sQ�6}�3��}�����TF�w11ʨ���$�0�t�O�5x��v3����!in�d��-��h�����s5�g�$A����2۟o�8U� D{?�?e� Ժ���eڦ)���c���gb{G��Uqc����_8G��,�׃���! ��������[��)�ӏ�=vјZ�0ʒu�>7H��X;틎�@����Ĺ�n�ԑ�o�����V/}���D��磑�wOsZ�(!������ͪ��w13�KM'b6���S�ަ&<�8�.�����F+�w˳ϐ����}�8��?�$1�g� m��ź�5�v�l��~�7A�K]�ܝOgf�^/*�ڇ�nq����آ��T�$�I���N����#X� ����� 2�ml��]�|�����}�NbΓ��u��9��>C�X\N�7�ڵL_/l[>I%i�k� �~�]�-Ԇ���kM�c�~̱��k�#=g� x[ɣ_U� Dk�����O�g�"g���M{e�^x���O�����h�ښcM��bs������y~�-�@�W.9� t>�sf�E����h:�A!�>6���ٻ��<k��g�"g���}���&� 5?̧Q��m�b��>�Sgv7o�w��q^}f>?��e��m��<3N�lLs�$\<��a;}��m�zT�����x M�E5y�:.Cxx�ޝ�o�%�q����bf�%� Խ����&~�� �ewg�����'M]��u�gE�]&���<��>%v��ޗ4idd�a�fׄ@��'�k��{�v�<�u�����}�ڭVh�u;��tl'`�8�q=�Ծ�����N%���'���"��`'r�h�;<�K�#Y�����*����]���-5ݐ��� rΊ"�^t��y����Q�9;�u4W�WӐ��V�>�r��ˋH�c�n� �sت�d��5�'d�����N��l���N��H;xھ�����&~�� �?�5���?��-� o����4����6����8�sϯ����q�4���,�J�"yuq��D�.�l|[�Ů�|ơ�r�X���}^(��io�dl����m�w����}���&~�� �?�5���=�J�V��ٷ*����q�>K������^�+��������2Nն��,�U{\ctQ��������;�b����o��9`�:'�޶B\�lwߟj�?�#�'��g����#�� ���)�e�{of�z|����k��z�QU:8��O�~�<�2���Lt�
�a#l�8K�<m?��6o�)�ֳ�'��4��仟���!�x���o�'̾����G� 13�S���l�Q��S��sg��u��)���r�wcALu��s� ���)��ԛ-��ʻ!A�"5��,�_����̓�n��J�Z6�H�;����Jb�����6۟hr_R� Dk?�?e� Խ���v�������ݛE[�i�1�Xj;!�o��w8�w����8�w'�d20�FV륖��f�{O%�%�O�8lvwK�2��M�>1N3�Q����w~ӷ1�֞\�� 2���#X���� �A�#�ߖ�g�����Ί����8Ĳ���v�<(��q��s���>K�g��jt�2�ٞ(%��q�����.a�\G>(��}�~�k;o��������o��� �S��ͿLD]���J�7�{Ar���E[ьoG��ގ�߫�l�f��d�/�F�6#���H�dqvp�l�|�J\]�t�I܎�͜�.��}���c�"g�������D�� ���-m�n�/Ns��U�����Ʀ�Dc�ϖ?��|sC)�lSm�%�ǲ�G��7>G	7�w��vv,j�3�+f#Ǿ��9�Y��ln�$t.i-�#��pW�� ���E�%?̼���� 0��/���_gr΢s�KԞ�m�ވ���f'������1n����8`u����=�[���q����=��,�Ɵ�L�����5��GH�����ð�v�|��O�c�"��S����c�"��_�K�[2�uޙ�^S�9q�e�EDE6t�M1��4�ӻ���B���R�{0�F>`# �� �e���}�߿=���t�v���5�Rس4,|�F5�-� ?*�d}��6������#�� ���/������mՙ�3�%ǫ�n��ѹF��zt�|�)�܆Wb���|��V5���\8e'n@�w�ޅ�#����E�y�d�ݎ�m�u[6-�ۋ������#Y��?e� Ԩ��A�h��nc�Z�j��9�l�sol��f����{�۶����T�#�f~� ���?��s1�%������I,���gv��n�n6���\��� fr8��f-��&)$i�n���=㹝�^>k���a����^�q���;5�l ＊��F���(� e� ԟ���Ɯ��I�f����4q�˚q�|�G��d�I �H:��� 6v��V����+f[-��Z���Iֳ���G���� ��?�5�������^� Dk;{�g����v�g���i�}Ү��{n�U�U�u��|u��d3��'�R�xDn���0uQ�;b�H�.��H13gn���>r�����y�~��?̟���D�>K� �M��l�S5Mٜ���[ح����(�E1=&<��=�!���[�m�/�� �=��g������z�E���оC��OK�x]ڬ��?�����;�vZ��[����8���d""�W�������]�lZ����~+�aޜ����,_P)�=�b�K�
E�{�H��vE����>�A���b�=�[���?�3c��qyS�,�^�w"��gs�,M?�����ybœ�4�Lva�^c���]��p�?O����G���nD�#�v���g@"N���p<^5Ѻ�ٝ1�~:�x>;��١�#ßR��播wH&(gbF��Oj�+܂�]d�x��x�pp���y!\��.����A�� c.iJC$��ՙ�c�=wP]ް�:�����u����#���X��r\ӕ��ː���咉�ׇ v�x����̯�PPp.�����Q�sj)+��<�N䲗f8�Gv=�%�la�I�6n7�]��d�bi��뻅����g}���Ϳ�^[@�	���v�>A�U�A���̫�l�ě�{���5Ŷ�^��wTG0�.m�v��n���X����ԲҸ�Cܐ�>K/�$񺔒nw,�G��爂W���Al� �9�O1H#pw�ܴ��y�Gʮ�|߀������.j,Wp�%��	�5۳}���`�{{{Zݢ>�I5?H}��ښ����>R�F�͒l���}i��s:��ݛ�._S����P���cqu ���kשZ0�፣f���   ; A�#���/AZV=M��Y1��{6�H�� .�;�#�;�w���۟�%��4E���ԇ��kB��\N���M{��H���8N�.���A�r���Zd����d��)���2u�q|/{�m1�@o�.��t�Z{e���f�$93�{�kn��l!�_Y�ŷ���%��TKb(�,����O;*i�zG�}c0m��~l~�mf�c�2�iገ���a�b�ԭ�?I�m�GR1E�-�=��и繭q�k��T ����v� ^7�x��nb�
�c�I8_�;}��|Gc�۱A�tvc+���%.;Q�p�����V�����&u�`�������;����&=X�WJ�	�R��)lB�����M� �΁�Gk�>%�۳}� ���K�Ǭ�k�m-e���,���u#��`=Qw�.{�x�Xi��.��.V��R֝�Vu���j9���\I�i��oj8���e�x��fN��	���.�L�Z͐Y˃������Ȗ;n�����-y�G���b8������r�R{�4��m�r~�۬��Le5^W_e]����b���U�ڕ��2�k��k[� p��.=�������5u\h��k�XO+���`o���;v��(>o�8N�.`D��ڱ�ķ!b�rD{�wc��G�#1��f4۶���t�t1��yzxZ��b��;�ű �>�|�7���ۗ5�=�/���� ��7�ֹ~�)?0����������kjDe����$������.����Cg�Ѻ�e������|2�p�\���9ka�X��8�߇~{*��o�A�_�2�W����ڞ,}|I6Y��;��UR׿����	<`6[f�Ӛ�-�b��/eam<^=�Z����2wGX@���v���e;��5 �Vx�՝��)�x{$c��s\9Aڮ��J�<tLi� ��c^��g_�oˬ��� �¹�
��ӹ�w���b�Y��6x��N�Nz�7�D�~�7}�g{�	�|�����5�N���Rɒ��C2�z���9��Xc�����-��oo\g𹩰u�����y�XS�2�m![s�׎�c��쾛{�\�� ��+8�5�u�z�GZ�?������.q�x�$�9(8N�����f������1��F�����Rl��5�o������q�8��*Բ֠�m�`:GW�����	����x��ʶ. ���Q��|�k�vk\@.�yPV�˚�elY�Һ1#L���)
��a2��17��c�z��Zu�Y��JƉ93w���^�1�]c:�7��[yvAsd�+"���lѹ�$9��f�w>%q��@��5�pA����e� �`�� �d�/Q��z�<�&�z�<�&�z�<�&��A��6�A��6�A�ɰ^�6M��y�M��y�M���� � �`�� �`�/Q��"6��@DD��_W��ص=k���Wz�	�9�{�X��R*;N{����/��" """ """ """ """ .7������싍�=�?�}`��.O��?��Β��ti�(2H�>�im+�����X�"�O>d��]ajn��>��`��O�3�/k����Me���^]��w��ƃ����-ѥJx�����9�;���8�#C��yw�=�(\g�Suꕯd2�����:��Y��k2֛^ؚx�j6��f��-��+��6�]���sw-#�$�8+'� ǿ�����d�'1�,ؐ@<M�=#��-C�=!�ґ�nV�ť�L���;o�;���o�oͶA���'��̆\R���۽�mc�튑�~]����p�$�����n	�AB�6�'���<gƬ^�S��Y��CY�e�٤2�A!���;f���ȬfjLK��7)M٘��l6"v1���-����Ϻ�x��;?�X����:�Lъ�N�	�[�󱳾7���k�f�o2�ȍ�#�p�q��J��b�?/��:��앚��1�0��p;5��ǒ�>��U�������R]�Ei������<�i;�в>���!�3�Ǽ2Va�Zl�\L�w��l'�pېV�-�C@��m�d����V������WD��trJz�K~	���u�B�d���\�n���Tѽ��� ����sof��4�Ӛ�����y)l?pln���V��A��Cw�Oh�.���d.����VZ>��6cK�#ſ%)OS*Ն�w7c�Ӳ�� ��#D����_�~[5'����A��q�r����g`��f�6��#o#����u.N�
՝eĺ����&�\�aؽ��#��j2Jإ�S��	c������+��DXܦ��)G6$n^�2�V�4�c� ��;s�Ga;��X�� ���X�� �[�V#�U����-N�2Y�� n� ��N��Pj!�2;�f�v^�猋(B��b0H�l�g`;r=��R�:�y)T�.�f�n�����[}����@�����ݛ˞���R�c!��_F��Z�+b�&��9� �+�q��2��,M������IkK�H� �>T���4��r�t�woS����U7#w��um-�n=�_=a��qg'�k�1�:����J2!�G�d�fؖ�V7��_{¾��S33֯V�r5��5��>6��1���,�T�� �R�O�:��m|��b���֍�f�X��I|��^Z��>N'���D�u�?���W;�����7&{�4RC����cy���m��{�D����Zn�}�V��0�F\�� 8�HHx��<�j������z9�j2��nkD�wt������)6e�1&-�o�l>���nqhw���r� �6b������a�ױo�h"Xl��r;:��&B�Sm��4^��	�}�� ��� �F�/�t��?9��p���┮!�wtuC�}�|.��n{������c�Q�^:���� �CYm 5��   �+s�(�����n�w�F�a��Z%��#��n�����ߵζ&���r�~��2ȥ�5��Cde�]iqr!�	�r-ۏ�!gbۭ5�Iy^�Φ������YQΦ�M!ۀ��l����\@��~� 5��[Տ��[-J�%l�g`�9���|�1�1��՚�����:Z��W}��*�cdk'�>L���q �ٳ�b�����LB�Y6g���#f|%� �xٳ��o1�R��DF�_)��V��-���M�ǿ%f�`6✗@�gM�[1��yY����>��M9=xKێ�2��g?�!�%W�lh�����Y��1M.���]�� �m۰���L��Wn��bh]��wRر�1Gj���t-����)�4�k��9M3N6[3�i�l�>�ٖ��c�k�VfM'slK�$}m����!�?K4n�aFݜ�|���9Vi�,�����f�&�t���uǾ��\!t#�� ##q�g��lԺ��t�֡�f,Z�:`p��]@�L�lZ%-X$�8�ۚ�}M��X�_)������EH��dN�'��8��y��z�M�~}�6�h�6ȅ��E�-����{�p�����t}��Ĕt�N��};g%g1�f�̎�D]���ї�oֆ�8�]���]�F��;t��כ/��B����S�䯮�����!��4�F�g�����]���\��{�ˑ܍��s=�dxv�-�F�5U�g����^����K$�GJ̗#lv�����Ø�t�����1�Y�vV�sO��n8�`��ؼG�n�=�V*k]?~�J�l�6�|c�����Q����va�;m�N"���h�u|�2�|�>��۩3e�V��״���g """ """ """ """ """ """ """ """ ""������]�lZ����~+�aޜ����,_P)�=�b�K�
E�{�H��vE����>�A�>��p��^f$��ֹS[�O���g1�$�́��񮂴�/J�_Q�;vS�r�˛5a^V���}�h��ϟ�$:cX�9�����ۦ�k,�cewf5{&q;8Ƿ�@�SAt�ڰO-�QfN�)��wL���ZԐ���q�Uup8�)�%���-��c�����V�D�����y�Z�]ֱ� c�����<�H noA��Ѯ�����7!oh�ZXhAf 6�}��o��z�{n�C�;H˨r�*�Z�k����<!�@X�!����esL�Fz��H*طQ��w�oԢH�'�62j���wY��%�p����;�r�j|N
�2�C!^����
pJ�;�$������HZ!�o�ʹO��v�Y��hO$��ۄ	��g?�ޢv*iƓ�
o � hIJyd�����^�����`r^������v��z,���b��Ǻ�ѾI��@���.#��+�R�GJdq7�u��%��-�k����G.�8�R7�n��Ҏ������7Z*W��vw��m�C�N��=�O`)͎��X���x�O������3������ ��m�p{�wi�<j?��~{�A�����ô�-'/'7�O�]-���E�3o�8,�~Q���Z����9ì-;�@��y��2a�c���'�(g����*1�v��������bݗZr�p��h,En�u����>*����Ù�q���H؃X8�%��;Ĭ�Hڽ'��'�>S�,��,1����p�I��H�� ��F����u���;��	�ӿ��>�i����6=���l�X讞j�F�j��2��4!��@���;����˙ߚ����pz��b��d�&�xb�^�&Nn�-=�ϴcͷb�öӉ=�!tu�{�v���ǳ'����>��Au�V��p��7� ��ߪ���mp�����Gj�U��xKY|�F�+Y��Z���0:�����py��Q�� 
ګ� �c?yqat�[:�i<����1Y�ۿF��d�k�"-�k]���. w������*3goQ�����,�3cռ�#����N^/�Y�܏$ ���=��jY����6�Po�M,��>g"���@���vqֆ���җ����������?��0�-�������l6[0��g��sC�#��n@߷m�;yӨ��~��]���lF��1K=�`�U��~.�Q��X��O�Ď� p����7,���W���&Q�K[--F�db�? ޶&T�$�鸙6/��;��C�޴��Y��&zl3e'!f[|\'�ns�ӿgk�H ��C�q�0�7�3d��f�Ǻ)$���]8��=��d�G0;	��gQ��X��ׂy@��$|cb1���xS[�^� �4���t�(]����#��N9��byr�Y]����
?�&��=%��Pc����V�tp�7��14�܍�&�r��~�䢧�X�5|�5ۚ���D�u���?���4r��� ����Y� �o�� C�[Qpld��7+	����Թ��Ҟ �KY�8g/}�����7obr��+��|�.68hL�$3>ȟ.:#��7m���|����k�ҋ%S*�96XȾ��/I#�� BXX�[��n�{�7��&L��ڮ��ج�#&��y�Oy�x��U���"���ˢ�A;�yH����Gg���k��[�6�+]E�e���u?yZ���;�s��+Ar�I&c,�1DO|���m�΂�f��,Mʰ�8���J�9��@$5�q���Z��Edtm[�ߵBӧ{\�B� =�u�����
܃���H8�LzG3��\��L�Y<#�0K���^>��n7bӻ7;�r��j+z��q�ז\��X�?|���w�gyn����\�:��-S����BkghY)��`n|�r�a���5�MJ�>ܤ0ѹ�����Do����p�����Ѷ�����4���c+����L��d�F̒L�l��^�����ݜ�a��TÃ�3��Ȍ�-IR�$O��ߺ'�^K�Cx�1��M�T�WH�������&>�clNɜgh�m��$����.t��hc1���T�}�3��'���	��N�b����#5si�d�L��9c�x��3����g{\��o���N;�}I6��fZ��1��(>Hڒֶ&���q�`-�$���]����L�:�q�p߸��� kǷ�~]þ�s�eg�>����Y���5lx�/co>���-�vp����r�fn��b����W�LX_Z'���p48���4��V��p�~�����Q��߁��ڄ�ɢ{C���!�RH�����������������������������������=k���Wz����|=_��XA7�=�b�K�
EGi�{ؿ����@DDD@DDD@DDD@DDD@DD����>�]�q�Ǹ��vE��t��v���Yj�j�N*¼�yz�\�4��nN��s[�԰�+i-G�g��3u�f .Ԍ;��o���]�#����o�z�vl|h�죠�l��޹�ż���-v��ud7��"�l���ُ�_����B��q`�$��FA��/��Z��=l|\No~�Ӹ$D�?�dnc�)�#��Q�O�q,�8�\=���ZgE���.��t%�Ql����jmÿh�6qv� k}�K{A�7�=+gR]�v*C��fa�,��C^|䷗�o2Բ�e��b���vk����,�}'@͠�f=�;�`v�n|K�gu�Lڧ_+��Bk�����n3��́��O�9T��u����R�M6_x������~���EڪJ��eZ�1�0ta�Gi���<���-�hp����I�/�PW����yX3u�Ǻ�Z�}�4r1��l�}�Ͼ;n��>���C%[=Fjl6Q���s�����yg��+OC#>v�To����f�G#��o��48,{�8L}�euj��d?�-h� ~�]�msrZ�p@9����u0�-��h- ���q�:�)�2��GԜ�8#���s�����4�z=�Sh�\����U�����s�3�㌴�yn�(-C���:^��^EQ�A-�f)"����GY��jCO�r]p��M�?���;��޶�[�pӭ$��equ���Q�P���xq<����9���٪t��ұw��˲���5'Y���6u�;��}�Ⱥ�\�[ϰ���3��a�0�ռ KO����dnj}a2zw��7��I�eiP������� ���vv�]%��3I�ښ�оվ����Ӆ�����c�����=�F�&��ӎ�����:sR�2�+�i	�kD�ג8�w�{�~%�Ua�4�Z�а����=��k!_�����Z�1��IRMpsAi�`�v!�*j�p��ƀ|G�� ���GOe��i�ܟ�nJZfa��b48�w@w>G�e�E��c-o��kE�G�G$/;���� �gn|wC��]>S9��b�:��ݚ�{������S�a����d�<��Ñ+��&�ٳ����9��q���%$�;��xC���p��}���f��~�׻�2�z�ՊR4�*��8�24�m�fd�w��~�aև���m��y��CX׳KuE����,���$��P{]�1�rh�s /���Rvv\@��#v�|<'�Ns��o���\6�~JCp��=�oK�le%l2囪h]�� _��ǳR�����b��v��ݭ��mq�nam9���hq}h�Di+\���O��c��W��7�����C��a��>�1�߶�ư��N�ޔt�~�Q
�)߂Ԅ��e�:��w��z��
6mK��?_	&B�r�!}����Ѵ�����?:�}�� �}KW蹥�iֹ�$Q�l|]�ڜ�֒{ �bb25��ש�&�b1$R����v<�w���nt�v�����2��N��D��!�VF�[�:3����ly �l�B��#_=z���-���g/� �*�X<`F9n�k��E}�^np���u�����Z�bN��!>>{-���٬C�.&iY����ī����O��쮛���`�j��gF� �҇@��cZ9�ߒb[���i&c,Nb����ݰ����cg1Q�0ױҐ#��qtm� �Aݮ��� ��Z�FP躥�(K��#^�>�M�A��;���nr^�4>w9��O���r�Gadt��Be.�y�f���sݭ��˽��g/�DQ���1>\f�8�$�k��;x�����򮧞�x-/f�|�R�	�;�N��6��.a�0O�n��c�kx�>?�m�g�n{v����}[n
y�4j\���և�!ͻ�$�Gq�A}�`������_[��f:���-ENjO��y����-�����k�v�'i;؋�H3�e��s[f�e1����<�ݾ-��I�N�7���(EK"\*���'gm�i�I�<��9��+��[�lQ?sqf�l�:ݙA�����"�v���Jt_�38��v��+T�KWș+fm��q�`9c`y����g�f�n�vR��9�b��6������۷n}��uޝ���ދ3NZx�L�d�����qk��������� ��}t��̶6��~�:�a�Wc��c����t��c�&:+��q]�.�Dw��b-��@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DD��_W��ص=k���Wz�	�9�{�X��R*;N{����/��" """ """ """ """ .7������싍�=�?�}`��-���u~���M���a����⟫��s9���ϗ5�-��Ԛ�.O�J[�C,a�׊-�;�i!l{	���n����>s9ѭM<�;�P������p4�ٝT���:=�8Hvn��j�/�e�[�
�+����=�����</i���$�9���m��B���[�Ðu�kU��do�f ��[�!������;�W��W�h�_��������A���ܖ:�G��O�w���y���i�tM��+�ܛ[s\����Oڃ�"h����IYO�G5�`.s�v �J��g��!�djd{q���@��7�'d禪ڇ9g���'�� ˖���#��iep%{vk���&�}�������%�J����ؗ3n\���@>��>�3���_��P���]Uk����y�r��U�H���A�F4�1�w��}��f��jܮ��bԹLS�.c�
л��^`�ԗpK�C��9�Ѧ����̈́���}��ˮ�<����r�Pű�y�:6�U�ϐ��Vr�f�l��G���H���CC�;�}��K����ӣ�^�5�HH�Ѱ�:V���ޒ��b�4�42R�ڷ�Qm9����ҙ]a�����6�Ⱈ�RHf��x�t��E� ���k�� ��.��� q
�"���Ǳ��p�pG���Nf�Z|�uÃ�Y5��nۼ5���8 �:L�� ��S���˸V-?#ZW��uw��{;$oi�;��>%�:?�za�g1�6MQ�s�|�k\��[���G�k��2u1p��-CR-��@��;5���_~�-N�8at���V�}�� �I�z$��)kL�B�'܋1��&|�J#�"ȁ�p��{ݼ{�����TiW���*k/�V�T���@��%cz���n{nˠau~QܿW��z�	�b�P�D�H#��9�o˴�)O}ېSa�t������>WѾ��f��2��C^ӟ/XK�����go�B�.���K\���������}N*�2}���yX��s3ϴ���{��8n��*����9ϥW)J�����:F����w ��v���B��O��g+��_�E����V��������Ku��a�k@;zN��xn��������v&�n�{c��ւI�h.; N��1���`���$t����񿼸��S���R����.6܌�Y+c}��k9�.!��;_� �W�ճ���c\.S�	�%�4�S f������,�lE�l��7J���lN��v��(>>�Ѷ��+��Yă�g�۵Rȼ�D�sY)��i<�Y�;��p��;})�LEɬ�O��'+�R9&�Vɉ�i�:�����n{��l.���#�TH�h.w��9�<Mp���!�A�#�<�Xl��j:p��2�An3�Ԑؑ�����V�߱�v�{��k[T��KPDȋ�b�gT�$�i���<Y��#�h o�j�Pk����\w�t���݉ĭ0���3b��8��nJZ<�	De��=��fi��߇n|��v�]�݈>~��g��b|��l�5UP_67���ӯe��z�K�Y�'!]�[i��L��Z0�CC����g"6<��Y�g1��mh�d���[3K��k���B�w#[Y�.X��v{i�xc�'�A�惩�ޛ�K��#��N*��ǟy���{IٹҦ���]�F��-O�?y:��yH�������2���6�\���7q�7�gYa��zj[�nr�y-CP1ĺ&�8�67� ����� �c��� ��N�=��j.������������5�V�M�0����7��P�7z]�����j\[b��t��$�YDo#���<L�ǃb6h�N�u>B-Ejl���C'���7�>g�T����w����]��Z�	��f�z�Yw1�+Z�]�h'r}
�����b���mQ�;:��D<���҃�\��?��UK��ka_��>:ͦK�U��5�ZKN����s�c讯C��?GyΗ��n�j��C�׍҇Wxs�6���q� Wj����k�j�j�k�I�V�bAps۰'�7XWu���г��̃�a|���nm��s���K3�k���:�P�u��F��Aݮ8s�<�պ0誇E���C�8m��?�q�S�75�ݽ�nsY���Y,ϒC�ց�I=�b�3���^�vB��0��U����<$샘���������X��Qe���:GL����R���s-����wcys�E���P^���� �Ϙ�.3͙�Ml�Mqf�\aǷ�����K�"i�r�\��Vk ���K(k �BƑ7 q�f�{U-�#N�T?O{#�Q���0�"��:���3����� �1t[�nT���Z��=}?V<Sl��� pY�Y\;ִ�>��ω����Cھ�'!b,%;���u91�ַr7D�8��sCG�xy��p�>�tm�-�9���0���fd�;�e��	Ʌ���I^\�EP�c�Sf�*^:'6	\�N�]cqy�40�v��O�}AGWV��l����gL��,��+��=�s6�w��ߒȷѦb
�&
�����J|mf��6xk��5�>&IVV��·�t��F�f��D��`���c�1��3(oVY��qp��eV3�M9����O)���[�<6Dl�����wn����#�+�dp�s��u��|�Z|�h���ZKK��#�#weo
#J�lf��x�A��.�2�b�N�c�%�F���8�A؀y�)tD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@Z����~+�am�S־��w� �Ӟ��%��"����_�b��H�""" """ """ """ ""�y�q��X.ȸ�c�s�G�;"�(i��+T�<�qV�2qV�:��D��xO. n�nv�-�hzw��'��m�5��*�B�b;8+բ���ial`	i�￳�rއ5V{AG��b�x��vT�{ϱ�M՞p3���4r�q�PT���W����U,���ݕ�Cq��PI��r��V��B9��1�Y��m<�;tYo�l��k]3��qn���n^��=�����~��/��|^|� ��pwU9��,�#s8�����A��^�z%�5��̄���Ӽ��Cö��LQ����l�{cc����r�v ,zYZy �R��}��@��;ק��A�K���x���9��Y��k�Q���l#�����X9N�rY��&������|�����Z{��-G@�狫kZLo�y����t�M���:�[9�̣�pP�����#c�� N�s��Ӱ��J�o+�r�R��r�qg����"�.��/	�c�x�%��!�����������n�f�<E}z�du{M�4��%q�̝i ?�n�/,�E�!�oԋ&g)Z�B��dmz��,r��2���6-g�WF��ϣ��\�Z�c��8���զi!�h�K�k�!��8<�i)s�}C��ϕ{)d���Nw=�i��qD�Ot����!Ӆ�F���ڰG {�\���̠tEy`���$O��e������1ǔn?2�c����c���p;�/3[-=��R�kM�ݶxk]��6pA�k�u~��Ya�g��f{Y��u��6n�;g;~{y{TgAg��7;�����kbe�s��$�65�1��$1��'�V��k�.�j�zL�4p3�H��� UK�5<P��-�Q�f@��ƃ��ލs����J�19����ä��#ck�|>ƹ�����
��".����ɿ4x��d�b��2`tl,k�C�$�f�{��Nv�����[��ƽ��v�9 i-?����6����bx�i�2�4|���v���z8�x,���{B�>�����I ������Ԗ2��O`���������=��C���Ϻ��+\���F��ƃ1F՗W��y�7~(���x۷p�5���}ΐz!��c���`�c���-���]񰸀Hn��	�~Em՘c��=�h�Q:�Y�z?ӗsڃ!3J7K=����7;5���`N��L��F�4��7���+:N�Ӻ'�	1��R��5���=��&���yTJz[1�f����R�O�nR:�gtY�=w0��<���\������[Y۸�w]8a�PG.L��� �� �,�'�2ƹ�iy�hqۈ���v�A�>?�l2�;5\S�d�֙6\K(������l��c<R��Xx}��l;���,��p���+�;�Q��:N��w{����	ߋ�nkf:a��N<-cw'r6�wzAY\@8��
�0Ff����N�2�*�nCTӝ�8�wR8����p�ĭf>��Y$�e�o��ɑ.H�6$�����׈�0�O`=� ��L �;�:�c=o�lu��[ng���s�����}�w
Q�*�-���xHx;�o÷�c��џc�SJZ�dIFKo՘��w8���ʕ%a<<���1��ܝ���,uz�%Q.�v�(�sv;�Y��J̏)NY�,��=��@\yoٿ�\�n
p�Y�d7�I��%^�Ӎ�ؖPm�.���e��?Lc袳�N�G��-���ژʗ��H��n���m����Gh�[E[��B%�<v"'n8���!E��xZ������r�y-�H\�Z�@�sp�r7���^Q������ѥy*�{��7C3)D��#K\ӷ0A�[3���������T�T.5�D�c/ٸA�e�^f.�ۨ�b��}�*U��������@:���u����l�嶓��+P��fq�v6�N���R)��[�=����#�nN~�8{y��j����������� ��=���L�鋎������z-[�}O�u^?7�ia�dz����->�x�5 tL�wY+͠m��s��tS��G�,3��[�u�Gjsd���D��Ę�F�!��{����A3Y� 	2<7c��s�V�S����F�F�6�ϭ����naNJ��8�K�Bx���k�wn�i�G�(]����/��pq2֭��B�o�u�K4p��${c��w=�`�����SȵΫjMo'dӱA��S��P�,͙�m��[p��zw�걙���X���Y�<\�Q�:!��5�t������/�����$�k�D\ ��ټ#�tMS�>��wh��_5'�~���$����Dl܁����@�u�zIӏկ�C#�]���a�E�`���2wŁ�A��ۚGCz��(���"=luH,H���By%/��0c2�V@;��cZ�7YV�X���Y�����y8'�F�I�B~8\L�V�%�k:�x�gb�t�k�yG1h:�Fٜ��5�wF8��;����ɥ���6�n#������]a��W��+�`itM��6GH#q�ŧ�N�E���X�FM-b���.�b�������Xי8�"[��[~�і������uL�f�$�&c��!���+�v�-;�H�Y�F�n��B#�ug\�F�\؁ ����"A=�CP�Hd��k���q`:��^fw�����ek�!��88���h��F�
h#��	r�e��q|N��@%���H�K|Q:gT�5�&,�&��RB[����c���|o�p<�\0��jz��������-OZ�z�ް�oN{����/���Ӟ��%��"���������������������=�?�}`�"�y�q��X �L����U������V�J��D於�Ip/�nkF���K;��x��4���f�V�^ Z\�_�y8A�Ӳlzԙ�%����Y�Sp�t���n����:F�[n;�S�lՔ�F������ �f8�N�\��:J�8;��6��Ǳf�D W|����[1.oWe�d��U.�-�d-v�x��ʯ���w��b��8�����Nb"���f�b�n�=~3�7G���6�g��<�k��hX�Ir]�ZI��J�;o���ǿo��[M�ԭ$�H�a���G��rI=���:�Ok6��{�d	]���=�\;oϷȃ�������#����Ӭ(����\��tW�4�s^7ydA�}�-�qW2]d�"I��F���1�rY*6���풣�k%��5�.��������n���ZkUa���d/��qI<l� �E�	#�qJ�)���Z���������[�XY7r�6�rc����d2VCnѿ$އDz�J�]�&�
Xz4�Ae�С4����1��n��;�n�*g�WCVK���˕�C��v���*6������d1�`Z�-�0��6i���F1z8�����Z�l�#����>�	��{S��/mtէ�b��-� �Xt���MU��aҴ{Q �g��7<8b0�(�EX#��ݮ�hn� �P!�j�$n`�.�0��q�!��Ki�<v`�h��c��A�Q�|�9�(�c���Y8���n<�< ֵ��rպ.��kY���ٞ�w!�u�6n�;g8���(,�G�������T`��Ȣ�b��G>&5�28LD����쑠� i��wR�4�vϘ���@w�[�Nݼ�@���r���f���g[V���&��o��o�����H�zrN�sz���5S���]~���5�u���#'`��@^�p�:T��S"(I&75�-A��4fX8# ~ĝ���ki�$i�g����9���^�x,1�F��ނNÈ�7�)��i�Y.g-G�}�,���nv.#}�E�Y��i�t�'3&���Y����.k@��#�.��͚{U��7/5�?Y����kxݿ���v� ��r���#�sA#f�F��F89�i�#�(L_H:c9���Ԙ��Z.��[�I<|'gqF��#��7��o����������c�>ˋcl�W|l. ��	u��a�0����@��=i,��;fchB��ux+�����֓�`۵l8H���@#ЃS�C#:P��:7���5�-<.!�� �F���-�ϝ+��6����r��nsv����q����`�ͻx�[5l�6�C�H,R�<�R�L��y�T��!d��գ%h�چ��K�Wd����s��w�=�O`(>O��)�����ɪ�����ŕ���}��F�&��>�H�+�;���v�ZR�Ig9�-N]Q�*�Vǻv�u�;w��m���t�e�'j<Kd���oD�$|e�qs=dr3o���T��Nޔ9b�Ե�d~7]��c+:�6���;�y��C�Hc�#�V�� c��u����������6^ ��b�v�3�A���'ria�*t��oe�`�ЖeVڹ}��5�G���ٮ�pv�p�+�=?e��w+g꺓��։K�\;;�c�v��v��Pq}�<�4��V̴���W��Ew�q����T�3	���>� �H~��v�T�Ѫ0Vq������!�b݈>�V=���ұ�k�7(�emA���y!���q 0;sސ���aR��?N㦿��V�P�n��ɛL��7s����ҍ��Fc�vK�s��+�;��`�6�]�fwIZ��F���a1�/Ac��#��Oۘ[�܍��w�qZ���\�,�8�Y�a�DH�M$n}�s���h�Y?��*�r!�;���-��p��[�`�oǏ��g��_��=�tR2�A�x ���A[9pde� 	Q�5��Q��c��[3'� ���G�蜠�]����^r��*W�;��b�G>HGV��.��aݝ�vi>��V�b�v:�YK']�H�s�Ⱥ������8D}���-��j�j�.�9�
o<GR��,�K'`�����!��u����w��u�b�����J7݃��r��O��>����Tq0�f��+.>;.��x�6�Ѵ=�l�v���1�'�.S�eؼFb�[�;l�[���F��cq&0ѳv��t쮱����d�x�sY ��ݸ�ya�4����m۰'�(ܗJ�G��c.j<e{�x��Y%��^�@9��`� ۴� �2x��Z�et|N��k������C�PT��LЕ��̔�!a�~�ө_�`y^��-��a�vm9�ڞ:�ac��i�����q� �*7Nk\��yp�nr(+�#�#'�8������h�(����۟
�A��-�]�Ѻ���s c���p�%���.�G���oc��qi�I��ȲwwXt��~����l]���� ���Wt���w����+�6e�XL��!��Yv���;o��ȫc�,�<�GI;$�SX�t$U���C�vq���6���0���an�|��a��� �V�Nt�By%.��X1��R]�@;�bX�7W��ܚ��O��T�ӿ^i��i���8|N&N�4��{��tZ�:�{x{Y oD"Y�9��e��u_;^%x!���l���撥���t�%�h��,QU{��IV�3�"���f�$lh9N��Y�VwE�lҸ�+�'s�;��(��?"町�RБ�ۋ��;��c����RȰ$��o�ܝ��� o����,� i��x��OV���nv{N���Qx>�0���ݱ��f\ᚣ���C%��������̂�F:g#��f,e�^�_'6JZ�e2�_�5�0���l7wܓ�n�D��v��=M����4��T�F�����a�p�Pjz��������-OZ�z�ް�oN{����/���Ӟ��%��"���������������������=�?�}`�"�y�q��X �T��[��Q��P����\W�M�c����ϐ�;<KkZN��VsS�pQQ�V���jk�$����&G�H��]Жo-�����ű��V��{���ɀ�8�L������Viߖ[�U���bj̹f�#�\��ц���E��6ݛ���v��!i�*ه�1���^�Aj[��R�������n{6>1��>�������3l��(� �G����"�ߑ� �t�k��Y`ys[#	�Ů ���8PZGDSѭ��v�V����m���x{|Jzň�W�y�d0D���#�ZƁ�$�@�P�g\��h�ݧ����` Jq�c�#'����m�=�5>��3��UF�xʎ���̱��Ǘ���;6s8ϱb�z$�Q��r�G��T��-�te�/�Z�W��v���<v��Gٲ�3����1�u�27��Z��Y:���t��^�\ys
5�,i�j�t���]�g�2�6;!�����Ż�A��-.�s���WrX��*T�Ҡ�b�@�Q�IZ�A;�!��<;�^KЦz8$�Z�8f2e`�ed�2���� 9�έ�����m�zk��Ěs�l5�^N�J�6Y�;�`|l#w�G4��9�|��]4i�����%ǲ~��(�H�`l�Ұ�H߳t~�>&��tu`d.�!���EӞ�CT�h_g�:X�۷:����ܶX&e�c�7���5�;�aQ�|�|���k��6MYx� �5��ϳg����CO��va��`�Y��gy���� G�#7��N�I8�C���2Lb䱾C-��:�G���?�7ķ<ޣ�骽ӗ����؞��B͇o79n�u��\��ty+��jSu����f��y�(5<N+�սUz,i�Q��]���1�m��\�${Z�������o�g��]#j�5���o�b��ؓ�̲��`��>�Y �ߟ�ۖ���4�H�cYd��.w�����[�Z�$Nn���w�q�f�����|>����2�qP�~/Yd-vݻ9rAѮ��Ct����Ը�Q�tт����rL?G�p���b�ilM������8��'8�y��Kc��v!d�=�D��5�;��|aA��D�����|n��d2��u�*ߊ[��\\6<��^�tl�"�Y�t�kԱ��\�EbPK"t�>0�2v���g��&0�-h� r��Z��Ɨ��s�I_F'�<�D�\�5��<-� �@*v)��nj��V"�/R[|/mi���㔴��}����&����F���M]��^�,ܤ�S)�'��qo1��qx�<�z�v��C��1�4��Ď p��d����'o�Ȳ�dj�}h�X�ٓ����4�'���}��c���I�0���QCP鹬�t9\�-fy#72�N�s�)#l��||'~C~�W�rVla���$X{��&>��q��������[g~Jq��NE,1�Pb�$�u1��c�q�>�.n�F�����T��<�8]��p��Ko����j�O���ϐ��<?�o�F��&o�n�޸2���)���9�'������GoW䛋��2Fې��N����V��2ǋ�-\��q��0��l�4���n��i�>�:fX\�q�H%.p�y��?�n�m��&�_c��T�1_��ɪ(gY7VzΦ�:�3?	ƻݿf������C��S��Kf��)�|������ⱪ�}={(�ml�2�I��ӊ�n��48��w=�����s9�v��K��_����KWfl13s��{��ۚm3���lch՚�Z�?���ؓs�8�I�ͺ����z�MjL�C��v�A����A�uG�R�O��x���e)f(�ł��"��8�H�yNG��&/SG��,��n��<��ߪc���~܁<�yB�PLs�#e��qRzZ�O��T�c⑻9�`��9�.������5�R�^���lщ �#q�۠�l謥^��jJ'j���*َ��Wl/��P�n;�/�;sh;�Z^S��_w.J��L�z�b��|�����~D3����e����B�G-F����W�e��e��mq��7�V�ܰ=Ց�3X��ƴ>�=�V��+w݃��s���Z��9o�`�C�ujѽ��=0�]��)��#��Y�n���v=��е>ۆV�k�_�w�nC�  ^��e5��d�X�{#x�εn8�^X^K�ؖ5���	�
3'Ҧ��e��ړV�Z>��R܍��9l�ny�H ��ٺ�!E�3ԑ�G�7>�F۵Ø<�Gb��z*����t�dm6w8�o�h�7��G>��.�+�i�n��U���;�@ܹ�<��%Fi�q�u�S˧����P86W�.G`FH��;x�j=#tk��Ykvq�*W�%�8{Ͷ��L��d|=��6<����s����*�v��͜��W5����IT�t`�P���~g��[���+	�n�S%$�i#3����a2�Z7 n|�B�(�>�d���$0:wB�\J"�L]n�<b>�m�s���V �r�[sX�q��L/=�f|�R�w�^��!�ב�i��1c�>�j�����d�411�"r�@;�� ;����V�S�-)og �6�"���$dӶ��+:(�������A�*.t��b�dvw�;-��GZGI]�d�|�x�O!�.�($�h ��
�SR���Ln��	:��o���(^�:3�il�/�T�ꘈ0uQ�ht=�?��gq�n�u�����ڛ��������'u}Sxw=f�$��;��F�z[�����-��p6ۄ�dk��ĆKv��qi ��d�+��t]���֬�zΟ����f��WC#/h<�%��|�uP�;V�u��jL4α��ӆ�I����e`{Zy��G"�Pjz��������-OZ�z�ް�oN{����/���Ӟ��%��"���������������������=�?�}`�"�y�q��X �R�i���S�s1�+q^��Nn�;�$s �ڹ���aڃYe�󴎡Ż��B�����#���� �Gy��dt��sZ-�L���|'+��>V�d������e������W���}�pߧk!ry+Gvj���ٽo <D��q3��]����Zr�o!��F���ئt��p��;�6�4�˽��ٺ�JzFf�s3�^ۯtpɸs��"��F������fګ,.s��X\ó�#m����m] ��r��1�u�M÷�߱N؝���i]�m/q�}���5�#V6gb��P��'ܞͷ��� �5�#s�|��8�U*۱��-�3c���r����q ����wz�euK[n�o��3����a�ٚ�	j:'o���bY��ڷnD��X������>���W(~�V��q5��2=�m�  �|-;����RiHhݎm>Kod%����!�c�z�8�A��� �(�7�Wۻw��:x�4z�'Q+hM$��7i��A��a�w5��j(��r��i�da�W�ٝ'SoJ��!���մlCx��j�1�;aobn\8��i!���Q�ŋ��{�Y�4HF�si'�5-t뇭��i��ŉ�->�b��I��a� 1�h<y;���fF�n/eX\�����4MI��uK��H�.Y�F^�8���8��n?1[-K1ݫ�^$�V	��摸?2��g[���������j8�o�C�/7�� �mc�F��3- ���+6l>)��\d���[����Ģ3�)k��v{ܘ��.�'{����Kx?�����"�����!X�20P6��@�O}3��"�4sq ��|J�kl3U�'!�Xcd��.-p%���w ��݈5\'���Ym���(dr.�Wf4�\�F��1�yk6ii<\}��Z����]_��0W1���$t9x�.���>����}��yn�'�>Zd�qv_-�U�T����6���9��H<�fGQk,&��Q���E֜�Wd��JZ�'�̐�I��	A�ю��Dty�t����cJ*��-�X�9o�nJ�>������C{%4�q�Cb۟�;��y�J{����^�+ڧf6��9�1�v��v����f��f3b������R���v<�@� �u���(�zZ��ַ����C4��F��|ms��.��[Ux�P���� �Β5��4V_Te+ܳ��֒��ч���c�@$Mi;�.ղ@�$a�ڸ7A�b�OI���⑵��c��i{��\@�Gw�q*��'Hd53���T��C�nR(m�͊�y�s�[��qͣ����m�S��\�Q�Zɗ���Θ��n��%���P�OB���-����$;��|����CJ�q�jȲ:�M��{�Sj��#Y�e����c�H�3{�G>��{��n䥱��U�GaΩ�mn����[�~.���o��A�_G�Dl4x˞݄���3�q>@%�Fy4����cK�CZ�A��t��֚W�6>�.�D��4�|��xy�v ���ŋ���-���6�U� �C_�Gq�b�[���埈�	�$d�K��/{;��FQ�Nr�:��y%|m`nw,�F�[���&iKO��g�=�:Fγ�.��2&��.|2��c�hA˴���cJIm�ۨ�d�X��,p������Mѓ��q�!�l� 9]�;��Pb�4� �]����9�~N�Ҟ��e�2���f�W�c�s�����cs^iu=��S���z^��[q���m�݀�Ni�t�-�k�j�mqx}Ɍ�s�qѵF�|���b��l�doP�[2qwDo�ó �!��H��܎���&�1���+�9��o' V���K�Ս�KN��2A��a�ZY�o%��O����r77)A0<g����ѭY��{>	�_�-sHoa�+fs�"s�v��/��O���ː�a�堍��ƃT���O�RS���~�J���g�!�WB�w�ڞ�w��Ҳ�es���.үXS�W�r �=�\�<��lͼD��-�]o'��x|�<E��0����5y�G;�����@'a�>E���t�sd�vn�_�������ó�=�4�;o��AϠ�9��s���á���R��lq�,SsF��?}�-ǋs���+�Y���τ��&d��i�y8�a<� �l|�n���t�CC/Z���ڂ7;w��l`e�69�J���Θ���cݐ�e����I����7��7���z�r����6L�F_�^����D�]WH�<um߶'pq7��b6-�ͫp��MfwpC�v���7'ą�=�q:���Z�BC^z��b{=�4��z9�j�����)�8k���Dd/�c��s�	�s~\��;����JkUF����,簻���k��ۄ \_Ź>-�ki֝(�tFB*�id/?���/��uøL��=��~[49܏-������y�2W�x�uWe�;��\�x����{��x|[���B���j���1�5��_�Z�畴'|���7i�H����ılt���ے�Wr�����.�7�0���8|;sq�b��i-�[�n��V1.?��`
o�������!���B��w�io	.
�߲N��ֺ�{/1ݚ�H+4�B:r��>p^ ������ևh6:�?���Q�b�c�o�;��]��Dw�ѧF�m3�e����u,=|F���Hb{�ּ8w�<C����w[)�����3ME�\궪����'����`��!k�zv�\�_��~V�s׆�x'�1-�f���H@������cp7A'Ж��чC�Gݱ��%,\� ߫��������bZH�o_�ھ���Kn�{4��a�lӸֶj�3n&?��n��ݮ �+`@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DD��_W��ص=k���Wz�	�9�{�X��R*;N{����/��" """ """ """ """ .7������싍�=�?�}`��-Z������3R�=՗�'���>(�Ɨl�^�H$�Cm�ki\�Mt�&�ֹ]8��1��O )w+is��|�<4��zxPk�z�\҇��8�.a������J_;��2�ȍ��Ρk��sQ�����<27-d*ي�b��V/5�lV8�l�q?���غ�='����٫�j4�Y|��wX7�9���Cw>N{�+��3KH�{��(<_{�X���\c y��o�v��'�� �����X��lF܈��(�9���v�*O~a.���B{Dm��^��R��j�M+�"���q� �QoY�usgv#�ð�ſzOf��L��2ڃ%1��`rIS����pquw��f��_��夀Fnk��ڣ\����T��guJ���o3V}w�y̎3�G�5���OJ�.?����6��Z�؄�\¶��	.�-��os�#`ƻ}������vo�C�a��8��ZgU��)�CD�c�fh��w�A�P�'/>��jZֳP�����e�A)$t}a��H�2��F�!�/,��8��������̄9k�ǹ�M������cp1�0�� a�o��!��_�3/Y��ZX)O]��z+.s+IC���pe�lx�R�O8z��7'1bi���hCF�Wpm����F��s��p� �X�|X�mJ0 �!��������X����a16�Q��I�:������a�f;�b�đJ��<v9�n̣0y��Vr�2'Dq��G��c��w� �A��4`��I捆���&:>#!�E�����N���Py��������Z�2�">銵Yn�`v��(��t}��:"��g�רunJ2��U��r��׼4�@܆��@��+O��H�1.��+LE[��sH����'Mg46[T^��sx����"+Q����}��9�3p8�g�T0yc�t�n�:\�2X{ ��6:�L{��y���~c��)M)�NZ���M�b�*˪ٌ��{CI#�;�7����i1\�2U���\�D��2�'��@��ă��"�	�pZuօ�c*GW�8�#m�w;z7*�3FQ��f��c$��q2�J�Ў#��'��y��[)jY2T��Rx�՞6��89�c�����A�Dc5�3��K)��<]evo����^"��-��2��M���q�bُ���|\|;�-���q��n�f��x�@�w�}��Ee�>Zs���4ta�e,cK�@�Mi;�.ձC'[^;5�f2�~�5BHKi١B��l���%���Hϝb���.���K����$ܝ)�W3�d��$a�.i�y'�Ų����ި��Nl��W��I��+� ��Oβ��)�f��QW����Y�;c4�|��7�o#J�q� cn��w3�ߝ��l��L�Q�66���sG��m�����{����[-��|\�^�(�.�����7'a�m��+���$ٛ�8���sz��ٟ�K�'���bCZ\OrO���?��lSXԴ%������|X�28�9]$Fv���\��,�o	X�߱��]�!���y�jkM�L' e�L����pH�aq.����N�O��1{7��N����n|��uM��zwg���L��>���z��;�dm��]#" y\�hV8x�hg�x�L2�u��tsjz:������*���̸U.��q��s�r��sx�i�}��n'U�$����?��lI�W+�n2���k �"�S�3�7�cs_���s�Z-썆U���I����(��k���i-Kqpu�Rٓs� �G9�y�ZF���}j��Y�k�Y�z�=�K��z�u]\�`1���@�����y�������ػqݨ��c�bGh�̷J��>��-;�8a�#M5j�7��Gqq?���㈷p�r����9��G��8���r#�*G���Z�9�Kas�cs��a���9�jM?����e�[3cqܴ���{Cfkt��K��R��kV�S�IӺH�|�oQ#dgV�%p%���<;ﾥ�~�����\��p¦B�68����)4��K�}�g.��5��z�������֯��Z ����M��a�'�+�"���B��&ˎ���i�}ŭ;8��#�A�b:̻R���;�3qf$e<{���c��#`t�#��y���7�FW_IVj�m�$��_n���x'���k[#K6 ;r;wi[n__i��29�u'mnd ���ҵ�|#�%G��kKc��<t�h]>j'OI��̑�n{�) M�L�VZ�9�d�,q��c�#nNi8;��=�*i������l�9�����������z}I�ؑ�A�=ݍh��t���覓���!!���I��q�A���nCX�]k�����z�s5R����rsp�!�g{]�#
�B�]Ԗ��-�N��2NŊ�X6d�`~�q������x���%?��U�hl�zvid/=ЛV_F&=���p���{O.�9ݧ�`H�z`÷VM���ؠ�WVva�R���:.>0�}�ho-���O��e��I{T�g?N<t����!�:2�Hz���ds̏�zF�Ϳ��'�OT��|�J���Q�e���'���1�9�1�^���ka��A`m�m�v71Vx�GV�OY���Zy���hyi�8��ݏ`T]�"t�<=;���Yrku ��>:*����p^ HCHaqwk�4E���%�����q�q���̗���o�a݇}�[-�@�6c�G{QW�v
u1��Q,mhkN'���!�_��ZX�{V�:^ÿXŀ���X��O�VD���\��|\\f2�io08��0=)b�mQ5Z��=w�l�%W	$���pc`��9�Ƕ�}�sA��gHc.�!z,�[%vL���0�� "68��5��\�[Z׺?��zH��{U�31y�|*����DSF� ;g�'ҶD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@Z����~+�am�S־��w� �Ӟ��%��"����_�b��H�""" """ """ """ ""�y�q��X.ȸ�c�s�G�;"�iiK8�E�s��le�B�a.d�74l�\	 �8{;|kj\�N��kL�ޖv>� 5���6��.��6���g�΃Z����'�6_9���9#����d���J��L�Q�(*� b��o�0����\�v�ͨb�)�Vo1�l3�7�Kwxp< ���]!�2i�zV���dZ�;bx�`�h�������K��8v$����EX���f��ۑ�1̭19�:	�ϸ�+�8{��n� kK���XLo,pm�Ø>q�(]+���&�ږ��D�{'��t��	�����՛�ZY��1���p0���٠O�ʅҺ���a��dX  ?��vi}�"x���۠��4��=�Y`GCy���Y���4����yk�6ū�:*��u�l�J����;ᆍ'Cjn��빓��C�!p��c�VOI�/���'��>6��[�K�=�<�(�c���3v���;>7�J��@ԺvZ1S��s�%��F%���S9̯�`��yX�tz�2��]�5�fk�����e�⊔��#+:���:Gq�����5y?A�n�U�Ӈ5r<�;/��E$wdc��Y��4����8���h���m�g��*d-R�>X̖��#���ل�7�O�=׶:t�*1��9�z[�[<a�c�����<�A{x@ۋ���ŉ�ӣ�MhY7��h �(-��B��}�],�4%��a�!�<۴��[�dh׷���6���p����?�9�Y�z���MM���ٌw�����M�Z�If�303؜B踌�X#�{�;�|�3��N�Ix�KK'[Z�x$.1��G#�έ��osy�F�c�z�	�M��	o=�Ղ��,�kK��26��!����`|���5-| �a�Y�d��N���[ּ0�"@;��H!q:{1��:��f�;���7��V��ێW��x2>P�0pn��<���{��V����M��I;�����G�Lr;��n�7Et���Yl�|W�q��u�����K^��n�m���)-U��z*J��I���U�
�ؒg1�ndMs��v��G:I�B`t묋��S��t��-�~�ލ�b4-6r|�73؛��+y{S�Gs��,o�f��Jc����S���r�ț<";�F8n�� �����ψ�̠����=���4�67s���~Ѻ])��t�і��l�(?;����X!3����w[q��}�B�k�����~�U�������@g5L��YZ���]��B���(�#ݻ� ���+h��X��6 ���5�f2�=#j+�ͩcB(�=�{h�G>p��F�75|x8��㲸<�r�$��?��5�i �w�8lv*^�x�ՙ\7P(խg��ߏ�t�m�[u?�,����`�b�޲+͔��T�Z����I/ ��Ȥv�a��v>t������;&fb�[oe��ה�jVB��#e�8�9��`��w'���&M%����:�����5�%�M��-�<^�6���t��n`�:�6�ű��ZG���1��	X^�8w�b	ޤ��F���49�� ���b�mABKx���G�sc�+�ӷ�&N ��o�l��c]ܬ��è���x�nY�D�M����+Y�n#�GJx	%�~�������/��P�yF2�*����gk�tҾ66(�a��08;���f�4e�����	疼,��Jǉ'�X�c�Z\_�!���������x��-2�U�l����i5��������x��w)w��m�۞���E��MFĶ��]�}+RV�lw�$nk���j�n��V�̌^?4,\6[L�Zagt������	܃�u�g3�t�2k��W�b�R��d�v�Ms����=���8�ѫ5����ۗs� 2W9�y��i��oe�������]�N��N�]3歷W�'i�g-'��F�t�ڒ���6��mw8����&��s1�϶�ĵl�Jp��k�.�ؚ�֩o$Ǵ2	�x&�v�۹�C����H�x�i����qZN�.��#�H����-���������o�M�r����7U����7�vވ�W�]K��S��֭��v��y���a{^�D��8rm�Z�G����{k7�B�F�B'����/"@�� o�r7])��j`�Z��[\��U�rƽŬt�68D�C�s�Gzy�*:n�t�i2��-ՌlR�bGV�G��S�8e�<�՗ly�j�ކ��j���n�۰g"�>:�]D3=1C�q?���H۟,�_EY-=�8ܵSg�l�֪9���sZ���f�w#��[{�]1���5���d�e�Y��Ӿ�lmllqq1F�r����F��M���t"u��=�T�Sbh�@���	�������6ߧ=i+3�:�#m���Z|��V��4�S�R�R�fps�O%b���&g��y�۩k���ў��C,t�D�_����\�� ��QZ[Z�5�6$Ʒ �B���~2�"I�D��7���'F_���;/6+����=S1}r���!��|�;����д����c)����䝏ȱ��X�p�x���%�pￏnJg\���������=3���^�
�C�8��c��&�08�t�F���Rjņ���?2緫Y��,��!���l�Z��|̔�=�K^|��b�GD��FW�[XK�����9�m�CU�c�U��-O\�|�\��(��3/��ag��,$�m탏5/_���t�4���9����9�0��wetU�;0�1�`�@���Vm}�4�ŋ��Bݺ����1��	�I$���{��n<�f��n�-OZX2�7LŒ�1�s�?t�Y�0	����c_�i<C�m�m:OF;L�-k�u�`j,�Y&�#��(ի�N�sX�~^�m�na�邥�U6t��d��Ẋ�E�O�,1��ش��}�D:�_�J��m��oV���b)��-������!���C���t��'�Y�F�ђ]'��=LQ����9�����߇}�;o�V䵽�٬h[����FܔnT������8rpش��v-���|=_��X[b������]�&���_�b��H��9�{�X��R(��������������������c�s�G��.7������ȵ��S����V��[�2��l.�2Ƹn�-�h�r�e�����1�bC]b���#6{\��X�\x�{6�n�".�>��##���m7�r�U��[dn7;�e$z=?�wO$�|�5�v�7#B;sf�=�o�8]a�����q2��R���d;�m�6'w<��D��0���]����;�p�գ,G�|Y�H��>(��%"76gB�1���ұ��Ӈ�iohA�Ov���E#K�NiTF��8-�ۄ�UŶr��a��vn���eJ��'W����l�f�I>`	*H�^�e��A������ڤy��x������҇Cp��m�I���c��J"��s"{���q������ɿm����j�SC'�ɛTq�Z�c���]-y+��@wx��`v�A�@V�H�Ѵ�E�v�ס��3��m*Lw�pq�l�����>`l�zf��u�ӂ�`fųۖ����.d]afҁ�ö�r�]��g5�Y&���J�����)$ �ry��D�ſ�d�����D���e����f8�eǵ��ɇv7����ƯQ�ҝ�m���d*��h٩BS[j+�s+����8�v潱ӥ8�G$X[�.��d�E��IQ��X$�l�9���G�Q���N�x �b��F�l?�&��Y�^�rX�1�2N�	�&�n�nm?2��n,�*��w��cp��p~b�p9ᛵ��@a�>�I~�{1�������̂�{HÜԺo3$Ύ\$��`$2���M������;�qZ��C�{^#�Y��@[�sߛ#��պ��Lf.��]{��pI<���9��\�84��	�a�"���*�{���cl��:S�������ሐ���PFW���cQ_��ǲ�;�����+#������c��3p��̑���9�u&7����3��C"n6~�#������m����Yz/�,6��������������>xcs��k�����l���nk?Vk��u&f.>����U���,�cK����	�;>$4&��Dh�>��wهU�Y3��6��y��� Na3Se�a������Z� ��wv��y�<V^�wS%����l�X��L�7 Z�|�T&�\>{?>�r��|f����c��D��ϳg�[���6���N��>��a�+�q���X���4N��Ȑ�5?:���w� n������L֨�B�F�*��g��iU#�� i<�٠Y_���
w��[��JH��j�"�엍��F|�ֻ�?n1᥆��>A�*v[�6Q���N9�.�|JF��5VS��5�Y3qo��:a��r۩�ߟ�e{-�q�K8���
�d�w6��M��/ �r�"����	��4ܭ���$�Y�Md��S�i���\6r7m؏a�xC�-�yn9uw��F���[0����[nvN�Wq�/w.�\$�>�\^5l���Xα��8���FbZ�s�f�cf�V�f��݈'x�F��=�5���*KW�>���QO5�5���Kܬh�*H��\?���~�ٱX�����i�����g2Բ]�+rH$��`�_�X����I�h����l�1Y�cq���ί3L�Y_F0��G��ųwR��b�֥�y���^&D��kē�,q1�-�/�V��, �v� pb��V#�~q���|4���ҭQ�o�imV�{wq]1���q���Պ�)v�f�5���ҵLGMZ/=��~q�o���%�gB�����=�=�'r-�Ϟ�U�X��7{�ք1R��d�v�Ms����`t�3Kc�E(q�Ë����Oi�j�����re=��
lչoؚD�W۪w��޳p;xg=�m5��j�cr�����.R������s1��϶�ĵܿJuq�؇��Z�U��agU^k����n����#K�x���qvp�/����j��#g�n���۰%E�l�Ժ{�����D]�Y�7�}�� 2k"�:�]G��>��x/�}v����[�NŎ�WF���Z���e)����X����Ӭؚ�V�qJ��אy7q�j���� ��TpV��r�8:����;��ֺC\"ap :B֝�>Gl	:^�PO��\�c8���̎�Qgi[�/ ;����;������gf�d`�Ǘ$WdL.e�����1v��������!�#��	���$�5�h瓎F��� ٷ�I��R�b~�!�1��QlV�i;�|퍭c\�ow!���y(��5隹}9A�޸s�:�9��lO` n�22w;v-���7k� �T����=y�c�'��摱�n��x=��1����C�mh�C��%H_�6����:��"��?`7;1����'Ģ4����XlK� �� d1�i��p��awgh�d��ᬲR[�+60Z�q��M�X�_��8���.C~N<�6ě�����g�!,�I�I�~ �8M��08��ۇ����;��Y�ۥ�/$jm��SL�n>�`k�u���.{����?ߍ'Lx����)�Y���~aŽ@��:�3m����m��!`����֢�k+Z<t8�5YJWI ,�K���}�;r�+~�h_�t5�귮A����"c�n;�� �6���G�o.k6�O�_�t���Ur�-|�Y��wetu�������X�V�}�ȱ��)j��ld)��u�c�0��v���<�����c�	Xz�[SCv����G��x{���p��p�����C}�J�Ή�Zf�-�Mڋ+[/ֆ4�,�W�|#�Czlq���m�2c~؅Ҵ�gu�s ��]\Xl{o�Ac��m�4�K�� ��arYe�+��\�#��=�;`Ii�\A��Oh}4��}�d.߹%�v��βW��� k@o�V�Ѿ���_G�gWcᖽ�6�N�S��29�l��q��v[2" """ """ """ """ """ """ """ """ -OZ�z�ް�ũ�_W��M��{ؿ����Q�s��/�}@�Pq�Ǹ��d\o1�9�#��kt����I��l6�]����>&B�,i�\9�F�l��in��nk^�Y%����p�/�;���΋�Y�r�q�ߗ���oM{��Gd4�:�k�����/v�&RGgb���-b�d�pگ�6/[�f,�.��d�CY���Z�.o�4�[szf��4�\�K�D6d� ��66?��f����N� ������SC=������3���Y���� ���H��'���b�-V�	Z�,{O��
Lh�&�l��c���2ˏ���T��w=y%,s�]�����}��}3����;���㺢�:���3�c�·q�/T��LV��%k�ո�����8�\�O}�� s9ф��VP��͎�>yi҂��@�k�]�Ix�Dr�a���N�!JkMq.��隃%�s9�}���2�-q��q<; ��6筎�����d���y�`��E���z*�X{:��L�V��n\͸v �ã�L�П�u�����T��Z�^*R>H8���qt��=��5,t;�_>k�l�!B�r	�#_?���Iv�sX�K�����v��t�����z�6�%3�� F'�kDb�H$5�v��g����ki��e���:'#���ӑ���'U�S���Y�2�[F,^>�8�x�`��k@��Bi]�m�I%��l��u�N���w��ͧ�ȵ8�ne�R�u�n^���+�@>;vk�b�<�Y4 ��p^	 �Ҭ��^Yĵ��0A��g�>�̺s�9���p�$2��?�Ĩ|�F��u�/P��T�E�ymz�6&[���w����!lZ?1.������drܬɞ�o����u�.��7WK��嬜�[Ew:8/V翰ջ�˱]-�Ѷ��;��"�]7���ws��{X�>��ݙ��v�n�k��Ψ��<�w[.�:�5nwP�����"cg��}�K&�J8̭,ݺ5/ۯ�l�s2�gDK^����H��4.�n�����1��s�.3��=�ܼ��o��I7B�.��sn<eX�g7��4m��%�'��76^�2*�)���s�w�ݧneD�zcӚwRY�]}�ڪ�M�++=���r��q�������s[}뢍9���D����=�ƏA	�N�gH��)-�R�;���}�7��6h]x28��̶c�k;x@��5���k�3q���7�p_��s�o��֝"I��~�L����91��&mg���@��K�\6����!���Z�����;T(������x۴l$gάk��`�$կvK�nN�`�E,$=��&��v��w䶽����n]C��jh��f��lS>0y��h��}�YZ��Lܲiܮzw�>�|v����V#hx�����ǖ�p���VJ��������W��s�����m�w���忍d�N�0zMٱ��H����˸ko �v��!�V1�)����6�`^�&�6ى�=��M����O�+0�M���X��*�d���*J����	-w6�;J�����������a̵<�#��\�Q,�o�@�2�nw��wܞ��uM#�vC d1c�8�a�Ie��c9�9� :�p�>b��j|�{q���[V�I4Uj�#�iY̴4���I�

4���GM�f*�:�u,�Zc�J�Fž��mPx�{�J�`�jd���fک.�q<�����Z�t�h�e���$��ǈ2�j��2��yArY���H���>��|yJ��]�_ɲ�~��G�<��M���9�quYN�\^"a${O2V����}[&Le�2՚�nc� ������~����Cc� ؎{캗T�MG݌��z�F��:�ݾ1���g�k�0��� ���o�"��&�s%�(����J#�mW�rǸ<.��rZ��j][����^���b�>&�%6��+c����^�4n��N���5�n]7�,�!����hd��)���qA>����Rb�ͨ��֭��=a+ed.�����c�����9[���a�Q�������Z�z0� l����R9�����7��y�y��;ը�|fbÅ��x�L�9G�p��Nᑭ��p#��d8ކ��RT��s��~�yw�c%�&�#h�$�/ܒwC�/�L������s�i�V+u��)��{v�l6;����1�+`�ۥL�UK����v�s%dƼ�Z�1D���n�� �H��ķ_�Ӌ!bfTy��y,M]�=�!�W� � �7hő�5[�k������#b^��xm�a�GE��:A'���̟*���s\�4�1��������܎�@6���Sz�>�?C��F����Q�����m�$���Me���l������ΠK��/�ٻ���ˇǓ�.�0��b+y�ϑ2i��ɒ~'� �����]���$���}�-���lk����8$o26p��ش}4~���@�NU�.5�~����u��i���'�m÷4pt?p�[ԳZ�Տ6�֊�ѕ������\^�!�q���f����b�]Mf�B�J�[���wTy	���7���Fy�C�U�:�1�74����6//���wetp��Վ��,y���E��Z�"���zV[Y*Pd������t'�տ���s���ѹ,�A6�a�`d�ɽ�x_fP����YXWi�gZ����%��� E�h���k*쬰���S�UV'9�k�'�仛���y鵇Q68��h�f0�M���/�,4x9��淏�#���.�'�j[zo�m�N��]f^�l�!���X��[� x ��n]h(�-��Ih�m��:W�O`c���������%wM�a��=/�N� ���G�(EV��Ɍ]��h�Acw/�ñ]Mg��=����4�����hsw#�$�jz��������-OZ�z�ް�oN{����/���Ӟ��%��"���������������������=�?�}`�"�y�q��X �]�IEO-�ru.ح{3L|�wPc���`sH�o�}��vl�%���s���+�\�S�|n�����ț+��F��8����Mx��K���M��,2�u1�n�&��G�;�\�l_c�����6��j��z�lu�{�\1�'p5�X��p����^��������4�NZ�2�](≢"8��a��Yn�ib�v��;��|�I�E#*�hY��zw�����4ف�����,{7iG�E��!�ҍ��\EKf �)Wl\dvo��O��2�2��42<x��ݮ�_����qm!%��� ��� �ۥ�M�b�e�ׂ8JQ,��� -g��v���d��Z����2��ߏ!T@�{��]���صv�3�f��b,���$�A�.gsW�%s]�Y������[����+(tæ�[�-ڷ��S�JY'`�Q�F�$!��nj;Jtӌ���~�_O �լ=B ����Ff����m{�w�iAP�b5r���,�O1�5H���#���#���l}�y�w�<[��k�j61U+G��V��]���u��i��Y&�=�i�0�݇	j�5V������V~�c\��㻜� �Is����0���->�*3�x.W|NB@��Ȏ&��v;��=b۫���z��b��FX*�j[S;���ll`ۋ��i ��߭0�ZV7�9��������zz�D���X[c���@ظ����ޞ~nK���j�᙭+��~WB�j�o�Ũ�H�l�dD���$�6M�w݈:��ρ�x�m��b�Xᓀ�� ��{KL��j��n9%u��5ᕎہ��������������6����Z�{2�k�WjK����������x���~Cu�7m�H4<D�q�7������������#��߇�Q��������W��Z�C�a����լΪ9sr6)"��68����m��+_�� ��������8fP���u��������� �K���H!Zѝ4[��I������Ø}'քQ�h#�c�;�� X n�r���`�-���O%k���d��2F�J~�.�o�N�vvmں�5�5%�jX�3$�V�5�<� �����\�ZQX�]�4wk:�l֑�@mHc�� -�x-�{vW��[T׵9����fX$a�2�d܍��#;��A5�Ҙm+��T�P��9N��;m�!�nT~��4�fcI�mM<Si���՛	2JjY�����x-<������pu��M���nT�z�����N^��@�Z��w�9�m��4�~�����cf���&�n���>-�I7څ���-�*�k%�d���q�$�{�gպZ���71Ż3�{��x�<׎F�8�eۇ�9o�Z�g�(�iMSwO��1���SS�Ԗ"��v���v�!-��е>�]��e0���߇�1�/��ĸ����K\��[��;�J/M�?��j<�v�J[�5w/�Ĺ��F�,f&J�u}`<sKC�G;�mM�rx{2Z��u,����d�wX�8����܋ ���-�Q�3O�P;m��[,����fFd|BM�K��\[�`>Dٝ-��8�c��Ŋ�9"�V�"ä���k�xGð-;�=�J�@4[_�:�5^���-�#|=u��H�'�����\�A`k������Z���W1x�%�>d���t�Y$h-v�C�n�wY�f�ſ%��B(�4�+U|͂67�� <-���Ph��l�M�l�Ej���\��Υ�� �@f�_X��y�dh;��lz7��f��M>��s{��ӵ����:����;� �7�a��W����~�+�S����5�^���m���=�y-�/vlv2Ś���M�V��]�h. I(1��C��3X�Yf�I��k�P�{H�e!x�A�ء�����f��� x�\��LST��Mj�i��30���,�6��,q�9�n� �����2s}*O�֮�7
la�X�N�S��]�6�Z�xO{�q;�m�6�d����@��Y+�c��"�ѲY���Q,̋���9�o7� �rS��cP�T*�	�|.oXv�q��i\�� d+iS�~���l��6h�6G亩�\��-K�$�p�\]� ���咟��[J����XQ��h�:A`��0�4<?s�@� �:�\��;RZ��dٜ��o.���o꺈$��o�7�u���G!ضm��k���ز��Q��n��/��`{C����Xx�l��cQU�Bkp���� f��$tQ����ā�H��(5���xbMI�v�fF<�sŕ��J�]����z�dn��'��¡�9`1ؼ�d��G�����Idc�!�Ź��x=�u�'pC[�}��ӝ6��z7�����l��p��[��k�i�n�o=�RW�l;7<����m;f��I�^�-tWejϐ���� � q���{Pf��b�������D/CV����%t`��nY��`�-���^��*e�ղux���p�Vqó���uc>�li��M1~��|B�!�d�m�	c��G>Oiߞ�b�11��X<|4q�!�N�z�c��h�9���z��Ֆ2�߻5	�>�������|=K���d��%�;��w��d��������Vl�b���Q������Ԑ�U�mis�I{\_�C˂�s�s�Y�W�k1Rs�oކX��we[d����H7݁���-�[�6A�_��-ڭ�az�(��K;��[ ��{^0D`���;o�`P�O��.k+q�ׂ�;3:.�u�Gk <���8����vD�~��Z8u^�a�ٞ�n�Y�l�p��� �����o�.�����b)c(� �JV� w�c�� �v^�""" """ """ """ """ """ """ """ ""������]�lZ����~+�aޜ����,_P)�=�b�K�
E�{�H��vE����>�A������յ��X�j���������#_����6��Ƕ�|\�At�����Qc�~)�1�nSe��Q' ys����}���>�0�C'�������Of<U�F4l���V���sK��e�֪��Y��Kzb���h�J��#G/H<]Lgp<�Xuzf����	�y[3�ژ�+�,u�6w��i`ٵ���� yA�߲*�]*2{���ux�H�]�*!�v��~6Hݙűi'�4�t!�R[���c����g����و-hy/p ����F�?���*U�R��*�+_��S����#��(�^���v��t�^��֘;U�B�7��������c�7�	v���� �}�p�.�q/�X�.'1Vfw����'�-����iG�o~�G=�z�+�˷-����C5��f���lvl�C�s^�7�?ڐ8�'�2���-�\U��%�j;�6�ݝbZ��s��@�#n{�s�pe�<�Pt��*�c�b���c�M�L���ۈ���f���[����r�$Ʒ�jY�4r5�h)CX���!к <]d�>"�s���_����n�앇�٧��V;o���ai`���y�V�������	2W�_aҙ#���0��SU{C8D/4���4 6X.�+[���;����ԣ�VI���hq �nx||��kw��W���܏wԎ�O~lm��y|fFlx�H��sϘ�o	�c��U���[`0�ꋸ���߈�n��ϴgC�mS7�7��&�1�j�!4S�q6�x@`ݡ�m�/r�"g�Ӆ]Gb<T8�_��tQH��Z =s\Ǝ	�q�ŷ3;��u==Vʱˎ���-�0�1�v̐��m;� �M�z�1��N�Z�ܿ�̓�}u�K�_��`f�hٽ�kmے�>�^�КS+�OO1C�z]\}��,������m�x�� ���z��E���W`e�%oc�{C�������5��ԭ�r�K5&���/�x���cf�"bi�r�b�:��EXO=�����Q��p2�+*�f>.8��f&�� �*�<�t3G:2ｔ�=��ź��F�]F~�2 fÉܝ˳�e�G�;T���ϝO��������������m��]�ߖ���s�!Ц?I�ۓ�rj�)r�ώ�e|Ih�65�nǋf���'���Fi:�#LQ�ԖY�Sik$��󻋹� �>E:�4X�-��U�Jx��^��mc&��/�98:�;�Cgl�e�a���8����F�ڂ��ێ�V��eh٢. �6b�����N��s��Ew�tt��9H$�N�,�:�����ix0�ɯ#f����XP���n����c�1=�&�xN���X�ox��ַv�6���t�A��.�!й'���U�.��`��ckx���#��N�u���Aؾ���J�Z��j����nd��v��ᑼ���w�%t�A��A����r�V�WAE��굱�+Q0������ ��v���h�岩io�����8ڲ1�;������i�������<�	�eg1�ELή����^I�ٵ�����4G��[�y5��;-�r�}��{߭k)��FHg��W9�n1��ٞa-h$�#������˒���d=���A����%6���}vVps:�����&�6��G1��(�Ii\~��؍=����X��Q���E7��h梴����5���Y>#/pd���i+��5�3��8�<o��sm��6A��B����f��Z�'T��O|��ы0�\�����[�h�׷r����1�ץ������	�iD�k�f,20���unn���WP��n�TF[$�OjH�jc��=�[,��;��t0�<�����bl�@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DD��_W��ص=k���Wz�	�9�{�X��R*;N{����/��" """ """ """ """ .7������싍�=�?�}`��(,N�������t���6.I+_��,�.{�H��ď"�T�ñ�����#��B��d&��6���X�C��%;yH�(�i�h�rdj�{x'���4Xot>�D�]���m�#��*a�Z뱵.G��#&s36;R�]t1���e�ۀ�w��,�:�G�;ػ�弮r���(�mNc	k�X�8�o-�" ��~��6���ԓ]��w9��r#`u.��ѱ����mNA�~� �J]�S����lnu�R�rS��b�g=썯�xc��	qc� �9�" �'�˪�W�ۑ;�?^���k6��ث\�gy���}Н �WٱV�*LM��־ȟ3e�p�û@�����Ű؝�d�e�r:OFQ�e'�i뗶6ñl1q� �ևp�f�p�}��*���]okU��Z�8b�%�����;7���@�7H.T���ʷq�lJ1O�Pl.Y	�+b5cߐ��Z�nv=o�����.K7��,���e}l�VK�2���Ľ�=�.%����1�Ж-�~,,Y��X��A%E�#G�p1��� ����l��%��h�[����4�f�w�%�W���=Ǚq?�<KD�Ӥ�޶�+R�5��@��̥*�H�{�[`��h�ȣ���ӱ;q�i�VI�Z��#%&�.��z��灷��ǚ���i_s��3�.��f����[!k�����cG�n���EО>"�odĘ��^��;L���(��ذ��v �h+l�]�e���n��VefXs`�?���1޹�����x���*eD�-��r�r�����]�.�(8ck8aa�O�qq�*��7Oa��n��Wg ����瓞������*I�=DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DD��_W��ص=k���Wz�	�9�{�X��R*;N{����/��" """ """ """ """ .7�����]�q�Ǹ��XA�$��c�}���OJE���7Gk-!�#$�4��;���ͻj귽�7�+�cQ�.V��jT05���L��Ǝ-�����N���{eX�\I�T��:}��{e�Mn���:i��{;����|�be5�Eym=��KpACc4{�I`��cKc��=�4���8�ȕ��΄d�N��V>���e���3�h���H#�����I�e�m���~mиW��S$�8��&���9����a�X��A���N�N*Cr9Kձ�qr}̎�q��}L�cg�[�]Y��Σ�oUo��㗯�묤�Z9�T��S-�����t�߻KIi;���v���e�fi��EwJ]��#%���F��;�&�X׹��`�-i�Gm�ŗ5Vn,V:�k�ʎ>ݞ�t�dmp�xg\����bڎb�e�E�]`��C�n���حGe�}s1Ī1�����&ݳ3f��zfq�����>��t��n}�_��`���<��T�ikI��la�n� �fkN���V�9	 �p�[������\r�W#� o�N���=g���&
U��kF�Q�CX��X��8�pZǱl]M�x��[�c����@4����;c�����R���듈�W����߱L�Vm������G��3V�O�oZ���$6,W���=���'<�8��c��kv �[o��?�����,�ʙ��uik�w	���ph�7�`Ѱ�1�bi]W6z䭚.�@��c�-/c_�]��A�r�v�ռ/���sr�� F?X�zl΢,�݈ϟ������v����#����O�}��[�b��VJ� \��c��˓ZA.'a�B���
�w5a��wS��N��������.���Ss��Un�]_��N��nj��Z������ <�A� �����Ϡ����D�Xg�w�_�2�c1�"�=��)ݞnk]��uu�A^�k9
�#d�C�Ω���$�����U�ٍ�jq5��0���n�z�V�>��������� 4O�}� O�'��>����g�7�О0,Ga�Ε��7��~w�\�]��R�������igk"k���6������� ��J�)��"������o�'mܮ�"ո��ϗ���}�� 4O�}��'��>����#G�ej�U�œ���k���h#�����`T��$��3M�8��Tn> {�>G�gzGetD\�U����nE���j���<�N~��?�D�Xg�w�O��,3�;�/��3��ڷ!Rih�V���+�N�H8x�ͷ ���~��q��Wpo�=�#3W׍�=�^�g�1�����gGft���?O'M��c�tZ���������?����?������2�<u�Z��b�s9������<�ֳgYޫzY�s��"1��;�. w���Gm���Ҿ�l�t�T�V'�� {?H�v����f��z��b9�B�����Ϡ����D�Xg�w�_���:���n�i*�+�f��������y���U\z�+1@�Ԥ����oz��-��w�mڳ����j��M�}�O� ����ϫ��@h����	���O�}�}l����^6���A�#q�c��#�y��I5�[���E-Y-C�ZK�ǵ��<����#���cgS��_��gO�hk�=������� 4O�}��'��>����SN���<Ϊ�T�<?���\�n�-�k�Z?�E^6B�)�|�eێ6���בp�U�m�M_�ON�[�F۵ޮ�������_����@h����	� 4O�v}��HYs�Z�� ��M �,B6�c=��%��ݼ�j���f�Z6��KX�� ��{�ۗ�W==�ٕܪ>?þ�n{Go�Ź�&~:�~�H�a�A��?����Ϡ��?����P؎��ح���� k|��o��w�h�scIs��Hӻ�$?v��G'lOnޅ�vcf��qg����} ���j�t�➽|������,3�;�'��?����)�ux;G��~�'�[k����}����'[U��"еO�����o�S���g� t�,P.�2�ZZtZ��z'1L����skl���Uq����DE澈DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DDD@DD��_W��ص=k���Wz�	�9�{�X��R*;N{����/��" """ """ """ """ .5��$ޑ���7��$ޑ�:�@�ќ�������>�f����_Ri�g{\6#�m�~�_�No�W���Y<6k4��Ւ�.�o���YZ].��ٻ������}��n�7��O�� �🤭>�QwIN�د���8H��+f���]�d�J�[������2���\���\L��4K'��"́�;���[����P�qU�k��qY�(� l��=�}��ݭV]�*�j�2Sh�	Zٞ��ىk7;�9�{�K�m��<� ��?l�&7���:|%���Í�,�A���qf��4���ۼy��m#C�F�;���"��>e�}���ڋ�-��s،�M �$��!y���_#�{C�3Q��n*�����_g{Wh�S���*�����#�,��CV��a��98�.`�:6�kk	<��Y���r�ڂ��Xqy2@���'r��	$�_��&����SO�/��WL�,S�/���_Eؘ�[\����嗢����'2ˤ5��t팆��xH���VCv[P`r-�M�ΎGx�`<�	�@�~�uM��:��Gkk��X��Z��k�r�mx�:GON�έA�>KR2�na���y:��s4$;m�ݛoڨDd�^��Y9&��hs�)��;��nA�	܃�~��M�17�Okk�w��g�(�1��n�mq�F#ϯ���~���[i��ｖ[�+]�H�nC���Q��~�T]Z<Fb6:N��5Ӊvۛ��#m���/Ѿ��07�'T� �������b>U��_E����?����􇣬�h���l�6���������Q�z�K'r�X�ؚ۞�d�cqpؐ���6�[/�Ψy̽��2U����lG/�4}Qo{w[W�u�����іW�{��s�pt���=���v�a�V2�_��d��Y'=��<�����ۈo�;��+�7}���X��'��&��c�V>���roF���������-섗}��lI`s�w�cK�m�k��
�e�A��e+���kd�Yc�y�vh����T� N�y��us� b>V���ʦ9u�'�O7�'���+N�q��d!Ƴ�w@̣߳�t;r|��� ,���uru}gY��x��ۯѮ���Kީ������)�1|�G�}\��:ʢj눏�����!s�e)0y�/���v�����.`��:*�@�[�.NN��F���^���	;���_��&�̂&�̩Ok*�1z~[W�iĪj�]_9�H� /�ftC��!R�0�x�� �0`���xw������,�BY,��+aoV���wS!���Fy{� 7�"�9����:��Uڹ���lG?�V��mî���W���?�����]�]7����26�e/���W�M� �n�7�?�WltK���3��Gkfu&h���xC���Oh��sO�G̝S|��S��(�|�}�ί�**�V��UU��g/��z,�M���~�XFa��%��{IXrt+<�{ƞ���L'ㅒ�����m��#ǹ�~�uM��y��̦{[UXΞ����(���uq�}#��:!�~�#ӗ�1`���d�0F�y� �̮S�#C#-��L�rH\�02^���w;���|�x�衉���S|��H�mq��?(��j���W9�<����������p�.囏�urqwē��G2}
���캣��ȓU�qm�c�[��Ȟ���7��o�|��0��p#��]��U��}|�S�[���錴wj�RG[�����Ϛ�ʆ�yr
��:�T�u�*�MS���fӲ4�4U�F3��""�{"" """ """ """ """ """ """ """ """ """ """ -OZ�z�ް�ũ�_W��M��{ؿ����Q�s��/�}@�Pq�ǹ'�X]�q�Ǹ��u��zs��~zg�����۵����"�0��k��0rv�����=�=K>�����������{���>'�}���U���[�3�>y��~v��L��>�ӹ�����N 紵���F��W��-��	��w Zb��o�62K6>"	��_�=K>���g�2����#��9��9~O���]���gz�fV�u�������v��Z�k U��}���h��ULS�#�?G��ħ`�'KMɯ5MY��������������������������������������������������������������������������������S־��w�-�jz�������zs��/�}@�TF>�B�՛5g��q�ې ���G�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A�����J��w�'�G�V��A���`� �O�X.����%_ջ���o��m@����s��#=���A�/9��WQ��v���'Q��v��� ���N~e�f?������f?�����%W�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�dȢz���P�:���P��(��1��_��N�1��_��A,�'��~;W�����~;W���K"��3���A�d�3���A�d�S֧��~+�aKu��j��� 2��i܆U�t� ݀��	����